library verilog;
use verilog.vl_types.all;
entity Trigger_tb is
end Trigger_tb;
