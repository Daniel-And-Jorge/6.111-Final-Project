`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DtbuQpcJqp26T+zectVGkmv5OK4mWShIpEVedtenQO4zrfts4wM74T3k9nKrxxt2W1tPWM0Wmnk1
Z8OCLhrM3g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d2i3th88eOgh94cMcBowDLISEdIQpnbxArCBVrpPX/HD4Zgsxjhba3lHOSbEcBQEOXI1mqJjQscR
sBrCpTdJP4j+/6ewEaQd7mINh2Z8/E3qYQ1sA3rw/B8unw8l+smmrHSMjvkG0HESDch2UYD6DiOd
DnzkOUhdr306BpIEWzA=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ILjvPSvbnKoV5EUyxxfwvyzjsMxc+lZdcOt0ULYWf2ZmnkElI+JyAfmZ566Cv5BybvIAbpkE4TAs
lbFdJpKI0wxt0RVWOuWLyVmxuNoSdo4QruYKvQVHEs1XVTIuysBzqE/vE45srqQBFh0chx3HuYsH
25NRSNvvSDfGVSbPt2Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DJLt4ZDDim1Hm/RC/uN3S28HGocmb+fp1NEHpBa1fctdY6Xa0dl9swUDB43bBqke6rH6S+aVFKvY
+VIXG+GN10oOrqBtTUlx2bph1/JtHXfdxrD/iDoM9kZAd44aYFcDDXx5Sf/dv44DWtk6Y6F1mpl8
JLJskCz/HtLXPFpjgPBR2FayX3lU5het3dp8+v5TVMXYmTNhbfbjiZapWjulNJHmNNgQh/0OXg9g
CVaGlzLERyylDYSPUDRiEjaCHzGk4TJIFiaR22AQL3bMyQcJgf9vV+5cq/llII6IkC1zQQzMnX0F
zMKS9e70V56XKvWAZvl54nsh7HNf4hYe1RK93w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dFBNohZIkCMhAoWOoktwYbWbF2tqJ762dUmpci7xJH+4DC2zZzFfQHC8adbAxdiNfNknj7dcVe2+
kEiX/hxC5LNOFwVUPriXwk4eC/0JE9Q0cKzIC42UDbXN7Gh+mUzPwxacEVqKG6pxmwgmw54Y+3qw
tPeM0v0WWchQeXuu8sLzfhAHySx759Rnmac039Bizpezjo6EzBHljszn7OSgYTMFlkPkF/xWBRbr
PtbvLsmJ77wKiJgiwrzsx00eSzHRPntQzHpul8zDvJ7GWVDjDYs1KxV+W+K5EbdA+VhVXdTfalgE
da0UFM277buLz6cWMHPipRcZ1BQpXoyLfH0Ntg==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M7cBjZ4oaFyC5MJnXQ2hoTYtu56oRbTi39VhEd3XwNgykupeLNWKfnTaF1F5XjkTEK+u7OKGP9b+
BPwvCCeyRMGToU3e6f+038OgCktGUmYR5K8IOq6/L1wdzi0fvinc2ZcnXygxPvS9CwChP6kQ+3nA
z3lVzCic6EARe4sKkUYVCLiIsTNc36CDJJnh3n7GyYLy7bhkSP481skgtiNmP7z/q+dfYYSqocgG
yETWD5QhiI2jRRuc3W3herl668378xA/1BlvNKK69Jlnh2n0iQg6i/b2AvKdgoCN0zpAv462oTKA
BO8Lpw0sSopNxXj/MEgPTpC3/+fRT4TdCtIYLA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57296)
`protect data_block
TkXIcuaIIkxkfSuRsCApwvKxVryahdwe+MBL8p5NKkYF9KpPLT37S8EVkKt2TeqqagnBDRWwVqjk
SnpJeGPk1SM0TpZ3fU8J0uB07776dmoag15+AOVYv/D5Pvz7xpnX34L34MZgkF6KvIyl0lbnC/fe
14HzUwYFFm1tzfz+YhVu8yfntWe6mgF3HcLd0+xh6M8+XgKJ+l4EJm5mc9KyaWSf7SdYWbVtEky+
4OPqMLYlyRGZ8De5oDiOCcSlL6wJK512UyBgAzgSZXW5f7V8at27AaemDrWUcWlY2sKQYFlDcow6
yoHY2yhZPpkzEJyn35pb0IE3LBtS37AEqT+6QA3CIV09LBoGePMRTSeID7ZHjzVs4/sMbCtuJY3q
49KcPwIH/dUMPSQZ25JXSKh/owXA8mkxeGBv4BEUUIuS1i2XeiPOSvFaam50RbVUqxlFWBqoovgR
E7f/X9lClQw4rCftWz+UxIXV+3t3OIvZYsMLHVxrJNeZQ3flKq94LXMUh172p57Nc4kN15+I5wV4
qvhP2JBAo1FFFIWD3eg5SStWH/qMsyqCwIZf0lCsVy4iLyT2Palzmi8YIaExhO1bOzMyassspmh3
kkT9SsyyNqfUjOM2euBnELr1dZwdXPdSNLSL4zDww6Z45qQizH0AMU8UAiqM5xQf1ucWIlLVlIW7
I1zGaatfZ2I5RrUqBAp/tLiITsznnjLwKt9WaF1iHQwWB4ghfR7Za6qqsrBkwKfNwRLQWiZFuRrs
+/qpB25/LXJqTA0+rr1WPZvOICo/wGtQLj1mHskBWJovNcAYEknM6wEZmKoomvc/m4usw0EMNx+2
rZH02j6Y1Dj08Ynn8OBSbsTYxyKsAxkhVPQUwH4F2+JIQlPKBlHhQhdnj5k4hY8dvT7vLr/+eg9b
n3IjNI/vQa9WLoFC7t4XtkxeChu0P2UmSA5L0ePA8RRQUmld6kuZn8L+Wez6Wj4vje7hFnLd59oP
hqOZ84YbdwyrPPsgzuh6dsPSkeInLEV+knzpiVNKVGdFM8OLZ/QYGakVDbMUx3GNbUCMUrrT+kgi
MC2iJw2lhHp5f0EaH3STQB2cdRwRqvL5EtuJJvZBvrh85IC0rVPJBaZs+6GH0hYQvu1Fq1pb7v89
VPJkwFnos6E0YcSW02mFZq36YRbZ/FbGjBIRrFXkaCB2DcF8XWQxwgqRqOvsnZJgoJ1N/VkloKi6
vNWrwpCArqlLb5JYpZaLK9N1l1knVEEO7n/TL4l7pLGwvQJtqJW/iEG5DNoqRe+Pv5CfU5GiCG/X
tLzKx+l7PwtUre+s1fK26g4396XBbXc5jV3hJEYzU4mC/akgERVJCN6YbTwM4QlBERTMojnII7Ki
bgULlO8yJ0bFrfhwU7orSpByLHQ2LHALwkKc7Ci3TOsgZ5/8IutFBl9/hdGsR+turBzjto/c8UcY
FOXtXgpy3BalOWr5OUnSajDArHs9kAhCy0NxJ+mKnYIpwr/gCadFvigOJjniQShHB0u4rhN2ccp/
zLXddNhg0k6UfgZgEZfKxavlUtEJ6KT6XG+Qb6GXsbCjkeej9B2wPBTtLZ+OtucS045CwjPdhrST
4HaTqp+yd0NB4iyQOo5hD85U2/Zqi3PCqPFLO+qlyhmd6Yk+ujPT4buHDXyl44ywTg5MJlbDwBPh
+IgLQZTlU1vNnRzqZ30yvwEMtkX6R9ECjdQSx/HrkWTAr+ddj7ATEQkQY3cz+4Xt1BnTvq9FcfvB
RhBsLmAy/aP4YX3gFMtGHl4bQrDkzy+GV1cApF5mqd8L13nV8dxeIS9Xp3Jr1Q+n3qq1BC23WcmK
WmjhgxdQkvD7Yyfb197+I2avBX8G447q+FRfbVyKa9P/Q7vxOVi7Eui7SOv0ifeI3lnfdEcTfucf
m0UvYQSr+As7yQ1y2b8MWYd44tO7YwosuR+GygnJNDvdf3s/4948vQpmyJ6x58h2D4DI+U62NBya
zaUrJziAEwv/6yxTeM4zJpO2/jGjwpjh/bYj5Mm/oE9pcxgXcOZTmp5cVm6S1GI1bjoGmSalOL5T
7CgVSPQ0GDM7Hwdu2AjdNevcP6UbMw0TwgXy+EuFGAGLBW/SHiLzaVY5TRUNFQRue7JZq+b2IPmY
8Gmsv7K5C00ZeoSs4MgBPI3QhJqWflUs4nHB85q6g1AKrHt3FmD00L1oaDwFa0G57m6F4ciG5Yy3
hrAQv3Cpptd8kHKdcBfJV3bEygXol9XChe1RXyGuDca+3q7of/orM9HMrnitxd0ZbyOkpH7HU+Zj
mF78gGI+ONXUBM1HsiyAYQaPvLfg69m76wcq0Hfu4Q/sZNOb34LK0c70SNfoJB4F8H8kh+RHSh2v
dsx9MZcFAmWnZ2HB3IQ/o/5uvdxW9RR/y6EVC57qD5QF03cjg+Y8YtYH38fN2JXogVICep+zaMPa
KQ3maAtYxx+vn/SCkt/pDtrzxUK9P+tFi3vaHIXevds8klPKY35vBBylPKLVUnXvBIqvFrLJ+FWz
X0ntv1SALEC7CUhq4LhS5lv1QFGgeqRkNLNG05ytkOP9irjc7v4rN5sBZgGtW13p8qmOLkSQXS3/
pqLBNjPnkbnV6HEmnxGPOzmk7YDR0SfqqbI6xTFV09EmX8FTDX/ZNGjFgMNwh6ePqWp4wY6ohHfi
YGBVtJy4qYVXWmlh5btF7rsD8mAsg8pRHXpbpF1xNWKKGcpYoacePcyRv//POf1/x1SGdGzgFScP
g6jeLXcaxfA89k25E2Pw8SR1fiYay513uxvoxtyvMlKiN6gc+JNtUhz2DBjWK6g0UmRIVJ4NwgQS
Qw+TFM3IQ9YtqHAJXcRrb3icI5TNd4eJmALGmOxBn13iTHMp2ocrEOXwIqrfwJMunWokZrAxrzEH
YbEbkIQVjur8Uux5Jt9o+xxHwrU6j9UswY44G+4DIncgc0RxDa5+mm4zzvfz1tNT8wNda0Ry06/K
MIv40FaagkmKEOuWzIUpbkBlNzd1qGBpT2xJnzPR3r9+pSps2wFa71k5lfxl+XP7hHIHn0+LjKJs
An7g1dgs3sFSbG3KP0JMevnfkW5oqQ3rnDtueqbA9nw6I87yiTu+3oKmrcJZkU6h3TmlGH1KzYs9
VFGsMlX9QbE1o7ZzfBZYFsOX6jnYCXgmJ1WyHMg3l7J4NKSxuKhxhqx7GBrl2vHSthq0BBhjDVK2
75iiAbcF05DPf/CFB5EtWttiW+8XtAxm2XTwHJ/M5/Che6i/EmWP3mOUvP1e3NlX/uIa8b3LaI7n
cFczmV3ZqdCXvV7j3YYVOXtP/CIzny26BLQEq0iQBgLSKVAtAE1s4+hRC7jEK96UGi1ObBtQDy9T
Yj/0wG1CvcpdHkGLAtyzvHepdu51GIzK44f8lToY9Az3EAsvWstFHTX7Zu+RHgye8QXe7YSkVf1g
YvJZNT5/yc45pfZttP/5Q/mz/NiOEGoPavgLyWDmWPLKcdApPBYGePVuyKDTjYUqtNQCOMLflzAS
PCnIV+KwGz1OYgCmRfea1gfKvJlCVJKMaUmVbuD4AAnRUQ2CR5kDI/x0ITB2FIh3gqCpTQkK3hAw
2FTGG2ghDXmzFVLWv6fed+r8M4q8EM1BmwkRJLOip2T2WEO/LHgIrqBIilj42vKTxdlJuqZ/stbp
ExavVodun4CuaVJdxkYNSx2flxBWjNtUx4wRhxT20HTkSgX+2E+Uoo8vKdtlr2LdQfRkfrfEueFg
ZdrTgQlUaR5kyShqqqlQV/FeFhQ1T7LNDughBYfDSigN4sae1v0WFhvpDzlJJkJ/dC495dyEzmu/
ODlgWTlBCQQ5w8xdHJqMZVuFTqaQtW0Nqa6B5FUUYK3tNvQTf99JJBSHTzpok5qQfQOcIW6u9A+d
f3NYMQ4ELQhp8wO59WijBdEHyVbGvQ0jeWuTDVKLaKN7T2rzMyV3bMEpSYepXg93mEOVxHghIYm/
3ZS7aon38UQa5qG3NC2wbyWM1GdQ1vONmo9pCE0Ct2h+SK08Y6HpJbzUkOXN8MqMhm/TD6Qrb/Z7
QhjgiE8tRHtSerJSgFlauJGPVCTAeH9L0NPw+b3lAzjM249h0xlDpy27ySGwI2+ayfsl2/Wgebdh
WjZBsvWsJgPsQBVNG1nG5txvZH18LSTv+4s0eCNX20MdIFfOsuuG68FsrOpwdBO1PZH9/JTC4Oyu
HShD0LFjJ1o8DFNwu8rIB0WFeerZk+PmCrPDVcI28QzPyxHXM6UNOXgE3US216NZ7Ex/yv+rXqVN
D7TH2FzfmowbB6uXqkhHQpAGxAjXgBMPePYcBkHRuQ2auzY2ysTrEMRR0jde0sDTlxk1+2LYr+AT
QJQqGnfz5aAhOcfC/mKqkxGgyFwLvm9sMcJm2rQauH7KC7iuuvJdlQAkIVD05Xkpk9tq6J5BRYsl
tJuSkhMnBEMT/N45+HxDaUpjziECkUz8IN+jbSnE7rRJiU/g4RQdukri9bel2W8vVKEomyy1Xseg
01QwyUh0VWobf0zcJr/SldjnFfxKdmdinSc8OaY0MDKnYH2La7/qedB4y0bMhSu1SCju6mj/a+LP
6u5KRro9a4YEu3aN4lhvikV8m1fQGDIbovmdvrZ/hVQUwuohgxoBnz9ayIb5Us4YEigPXvoX95LR
OhuzbqZaG7To1tyR83rCXL/EaBSYddns61uW+YXc4A8O3B/bLWKaEQbCtLv7kAKfXE4aRotCh7uK
mFEmNKsn4wvNziiNvZtS0jEjMTHmLvTHFSh/jLer2JdTWD+ICL4sksgJQzbov1HsNJxoGImrpQRX
aVkJObMSAr2334aTwVv6/shXsgvb1Ra+HY4e5a2DdE0AHQ81mfnNOJ5aWoaTtTvuH/yHulTm/vFs
l3ngaBJ3WCjuZAmVTkZlOC1Xrcv14aAyM8DiIxPjDKptbH5Fq4dRfjVqy0Idj1BsKZMuFWA6DJHn
pr0fUEGrEwKfiLxJiOOtSR5MduT78SQRMbxmuVDqHXZhXoCeRDxsTxnQLG03+KHWHycgZbofcdbE
I8pkt5SXM3buxaCL6AzCdoY7SKj8HYTklGCxPeaAoYSRO+3raWos7MP2BP/RuqMbMxFgvIonSI2k
zGu6DyopQ0BAdl7fJRi5zx9+7b00SokhUucCflZ52kfMg3mLQa/3E7wOg4DUD/Prs/kAzKBQjkgm
kif+vVZx62QJcHbXmyBlehLlUcDDyZtKII5S5uc2ABfAaaoDjrUvcB0gMrIcYam8p7xVcm1TVMxa
XrZLfktbp11kYSw0BMya7Rjt0MN9dqRs5t2WRGNvayigO5w3m1Wq4Zeq+DQIxKkU3EKi7f59BWor
eUvvEjaewFqP0rkm3L1bV9+A1apsxXq/Yu08eD50HxkMt7ou+GbPrbt6sr2uMICfZqCMTDyW5SQY
WU+wtC7/oIV47Wy0uC1nwIswqoDtVyceuAlfwDGvDwSokE7d5DJ3mhwS4CKHJc5Q0rzvFZFtoH90
4k45X98dtYU1Eq34ehAHpAAqSgUtn3M5WsgioGQ8Eg6t8Oaq+HC+AxQV3eCajJSKc0j4ogPbFpKa
wFOyX8BFngzWgudnK9PAuKxQOFXofp6rt0hOAcsRNzgEdY8upscA/fBezNJHudxFYdWMC1vdlx0X
BgqrLH9v2pqRcMgCAIfM4cVloZxhhYnWK/EKIcnQgB8nhsifncf5kuwasmI8o5fKhf0OrIC2tCRM
+GRlFlTEUtgTyEXaJppuC2UA678xtD7J7iabyEwSlq1IjXmO2MhizVuuRjZtg54wr9koyQOkZM5o
1D+rbJPL8kOBUF9x5j7xNbSucu3s3gv8FPJ4MSkU/kJbtRNuLMSLFwPNZZ9U+IF6/L0O3Ap1vYRx
hsT2/GCQ+B2jN8brLmMIIa8QQYd+GS/Mq7k9WQdzgvyOrGDT/DOK4s/Dv3c5Zp2kcyxG/EfatJSm
IokxIEmSEy9Af+GLIYtKtSGtruBE+CrJGsynK8PDYiXlF9j84uXr2Yl22wf3X368zNFhLDV2WYaf
BYMON3HvgNnY0l9rubYOC1Cj0OVnN/YJCzukQa6frS2BCwukFzxFtEx7YVg/iFbUPdkSmOuFBfoD
B+cH6UPPU2ZNjmfL2gcZpXhRL4szS7SRVzCzt0lr/4O4+5YrJwEnnu+XkUJfTtAK1N966N9Yk4fG
YZc47GvrHdmVbvJygEvPmMD7ZBWoHA8RSVImXhQknxnSK8XzeQQhuJp+D2+n+vhBsPLx1ZLbB2iw
hPWylksPTR2tQgAfcLRpuTF/96wj6wqKOEIA+ZbxieX+DfRwMXpeK0BsggZn+ZKNvUItfNepyQ8j
z1AI6tFXT7m9K7DDlJ6AOYy5XYDYcNrkB4gU36AqnG6kKunViNJkV3Yqjw2RUS/jjxrKiMcBzAd0
HiiPQr9O1DOoeJnZYycDM/J/QUBsU+kUydUOJo/uWk1O1yvbVAXquJ1u+h97pLjBYE/gZ5Cl39Xf
7b0zgTn4etbKw6prjM57iA2PA3axsFElrdAos8lw3IEceJKiNALb4SzSB1yF1o2eAspOS2q2qIa2
dPeDTgEuteUXbwLUC4Wc72xeRM93sC9d6ZQS5CwLBj8B/lWAesP/qh8wBQzO5NJ+lt4qEOUN15Y8
+MEOqHyafq1jxiNpYF6pEhnEPzDuTchVJgQF34c0VXOqAIjn/k8Fd65cimcBt1lSXMH/og9CarwG
9dmgZ4UfNni6jtGFdfRPmvpBG1hDlV6W4Ty02kclwEM0iwYXVkp4+VKu1iEEYv9pMLQ+FCK/rEPQ
d11Zsg6j9Wj+OBS4zuNFLW4Yep+Wpb6VySPSrNMHxMxGIJYtAPTNot23FoPKPODGN0vYyQbfEwVm
uAImaGJssHUBlgb0KW1trRLCEVmF7nHK8OdFy+EiCLea1vpIUE8xKhL2k41c9mRLS2YcLz3WISeO
KNlFwNaRQ+hLvnW63Knv6ZVcphneMh4v6UwwYJU9RmBFtvBBVLqSHyRhkYzxW6bwXojfCY4NGjWY
uEgJsH/7yuP/Xulp56VieuyJavQW9iCn9yLGX2HSR2OpLc/Q2GCQgaMTcG1dz1rri0/noZ+whelQ
NG4FvnrxsmWF8+LLA31r8bslrwwdjEsKB6vgmeFbxCsPbyv2nQBNN2xhHJBv1ntQWHMulSKXHz+d
2NkOwzSe+p9v8UGVi1k8deGgPs7BnKxZQFIrq+f9Kc3SJ4X4n7cUKwr4b7wZTGdhW5CZdsBkvssi
qfNZyDnwlS9xw8ncNWdkllJVqMre7CsHfdDSzQIJZngAmhmfOepATRKd9S/k6M2oYe1DEBMmNcZC
jnngayaugREN2axLZhr6ZKGP0VkogsAEB1bwv9JAb7vlGf+XiUthlmVbudC9FkS3yj5R5tahHrrf
UAr6v0cHK3KqPlXhIeoaj8MX5hGkDcefV1kamGNsicPbpu9IzVOwu/cWnTFzRr+Ctgj8ntkhaRqP
SIqlq7ES8wL/6WKbKizZylj4bJ+9rij8oqruBTgfXTNvi57hVzUkYgB9s4DSSy8lhmq5d+htEMmg
xNiQDJ28hCCqi/XNoj60qrZAJo2Q1gsbK1yUF6ZA1qDCUMyhAKC0AfACeLe7jP1zD3bNLNY+XAwM
8IutaCcaXyvB4UCuiDV3Dpm5a++Qvc8ReOJluFaNFV/rYzFYMgIQnK0I50FbkjkW4cJhGSEYz3XF
6jH/HNkiDB8sEIq9EWqZBu1Iyzur9zLjynazZIrRkAzOSdmLsuhiClb+Odq7Hs6Fc0k3zUxZ+I/U
9+PSuVxSliugwMvZRWsatcmU8HVmAadUEH/30zvKxTbhaG0TlK7koAtyxojfwMI/OohbLZqg72C1
M2Yofl9vlSxObBA/XOJMmiKKboGaJ6Y0Sl/ceqFNPiKYdaPVZ1q7Oqc9+kF01ZP1OL/oJSScH1dZ
Wk/Mc+MQKC5BxRBe7i5x4fti0otD87xlj9B0k0JVXLJyoLSVNM9AySNiSKwrj+vxJANZ1XXw8VTE
fHJCQz9cRlfJOzV5YjTDyoVKl79B+7YjvqSd3zBmBLbypDh4/mjUPf2W09E11UdDW5uMUKlhhxrs
1SR8zHSxouq8idTgfJeomFeptUlLx4xdVlRXzUt8yBRkXd6REPC4YMwrCfgLsUl8Bw0YG2WbaPfu
XlAGwJwP7BuwotuZpIjGcSwkwDKemBrVCOZfI0W/EpaVVs8txLlNMLVkNXNpQE34eBLr+PFhn24h
nm3GfH5axVpjAN5lU8uynz/G/4ckUS3NGBQJX1sd68dvRJ1rvK3F2iQ+lguJ9lpl+NMDKa+sL86N
zXFTQ4Renv03CBfqAmHSFgsA+jjYjQ5kwXOmH7ipV54i3mf7DTIBLs+zh7bI1mqx4whU/A56afZ/
ax4i3Pq3M0hMXBa5tKnYCjrIXCFtY9E0CyLNJrGo0QplqyaJjB369ECzmtHt2GtlaqJHbtAoDmY7
40JEG+Kc/s8AcHKU/Ww7IrUMmWIyNqKQe+LNnYrPZmQdc+ARJ1pUt/TCdNF72D8jNv6AutfRxvF9
vxa0ow23NK9CxZtPpzmef/EJKidstZ1OzhJQSxgqTbu44XhFtE+Nv9qaYdYW6m/SHEYEtQT8R6tB
XyBKKaOfNWS6y13PCNnfJPGM1ig7TNOm1fREPrV5eiVhez6zY4Cljsi8tWJusi4Q27SPgDZnmi/O
zYOgQDtDUVlI7khs5aiovfLUImEiLMm6xTU0dE3YVhI17kV1UQYiUR7bjeU5bndNanFNRnAZihfV
S24o3v2RgYQXxwGIPjeEhL8QjiUi6ax2UNjNQzopyH9GOIDKovh/WGtN7z9d2P4L1igxAdwm9BM9
lHc1m/11JolOJ4y8hcEtD7dO89VggzfnPRCpysjVGJs0RPXsPs3wgvvuiLJiiyXB+JquVsEDcCTM
Dl+VDmrCB86Xi7LERnnwhDgSi6+38YFMfHqDcmAwIaRtPjMRn3qglKp8TXtKpRJl5/V5jcJSgOgl
ClS0wt7rLjAYkixffnYwC8lq4zfr6S2xZLZAOS1aMgFr5wg2hqdms2n/TvNJgv9SuHlBHe5U2XIB
WUSY4PBmi0WZ2I4V31KD7wWj13Wb/Ucab2/46YNbHR/fpjCNs+OXAZRr/aVaz4lMZ3zJheF67Ws9
qw/0u5S86fXAPsiHZwcOCkUlOxEZm7t7dkt3cUTLsDfJ2rmLqBW65lTRZzoNHbHxxoJZgji1kj4r
MKL1+raUybRcMFMBWqYv3V7FQq4tNlbk2ZvOdSgktJytLoEl5khz8NwqN3lKe9IxNa9gUq2xJQ+P
HEQ7hqgVCIWD67D8o51rse7Z6AbnVIOfVvjPuCEQn6HS7zl5we/b+W45OXwN8PcQNU32CkCv3uDe
lsqvN94pSyPlmFeyrzK1NRFjbtt7rdpSiHKruQIZ5DwAz5np9uMimiQYr6hl6ClBP5ye7cqbmJG6
QnryUkg2oWTHbXJ5IimLsfVDw+sHVjje4LD3PgB/JOu2yhR823/JNSzK11j2CTD+tuEjdYWAqaAS
Y9cwTBfw//6BvHpWBg9ioYdy8jh5Q5zpC0OGygq8Y0pwspHVsU4Xt7yAYQKisrWZ62vBkrS3QjvQ
tJO8iEsDV8QGFT3EPPS2uk8axOaKRJEnkYKcMhpwargqzP6sU4LPZUUTbvukIikSqym5S1v4JHuf
f5sWGgphxN8EkcPBEO8Tcj677GK4SX5NMKh6xFRopS/411ARhN3urk48n+EpcMiC7mEvPon25hMs
pENcRieMmATMXXHKJoZofvywqbl46kmFsxqcJuuEsg+gw1xtOWPWUNooQoOK9SsSIA+dIs6HPrpE
IH7lP4JUOJ8Uyp5hRfzeWwQ12QVTZGUmssITD4mEMm1jyUo/0KpsjCwN0LLge+CF+0N/wSwFsE39
XF31ybnz8bbJR3OGQJjw0iMUQw0GeA4sZeWR9VL2tqkfyPUmD++jtyHoYXEQyqQE9GnUnLViEYTF
jykQCIILamWiZaRqk2lUQIdNcO8h26pupt731AIQbKhRiqh20j1Q3pl4LpWlaMCc/D0rdYQbxoLJ
rYTTl4+ET3QgqCjXNGySKS92WSe7iVnRSaK9vQs4QC/JgeISQO3CdFjzDBKSs8folpqbT1DisBJz
EDbBayPxbUVfWckXwShPqCZ8U0giFpHYMfNH/Np+JIM6757kyLM3SvhFqXuXh0dYvqWLPRfC2bjg
boZwAD3F0rsVdkKiz2u5b5JCLA88u94HOHPoZkwkj2myOjj9uOcdaWSkgazOXhywQyYAFK687EEB
SYlv/9UVw9ZFFvebOHc+sVs60+CWXTV+v/uTBeVckcNTmhek9HT1jcfAVwqZsPMuyTNEXaenzXUp
RzjJQnn0rcNIEU4vPEXgCwAA7NjhuZ5pphn8jzVYPyxe26usGo0racnj2q+vlh38ulI/vDyk67Ea
VOBTr92KzPdS2uhbAiChur8R8VqZ437HVs23fCBRd0jUgS+SzZCVv+jUenbhgZ3nkdAEkOqmfAax
HcYxFvm8uGtdHg/URABZtXPIUbUW5cAHY4bBEhsmS/bu+KiD/asIG8Qc58w8vqXygDE2NQyefwXe
y+ntcgX9hSUGh0YX5DIoDPllXG1EmDeI72eFXx2T3aRaQdz0B2YoShF4mSr5xBy9r+0mFReiR2Un
FOpvZzVAs2hl2fctHjFSWueaIea83B+TEQVMDExey4c0UsnkwMg6bz4WJi5odEklNtxbvGGOUXOI
Z9bMAjZCL4ae3yz3sFdkh/fguEqi5nfq/M5R++ZVUiTTV32mNr8OTRMwYm/P1/88f99PA43dG/FC
QT/OllRY130chWCUzZCKP9d1k6zwiLASdaigaNtspXzTqVVMgAizUAiboX4V/EFFVG4X1SDoDR+s
20Z9xgo17JdTFes+xjsKGfL5wPA3YjUzeuYrXuxo6Fi7c24Vam4HWN+zZ2LznmdLT6fxtHZhAMy7
XM1E0MSfOJWaQSmCmin/f/WGjQLIWAIHntVS1yiFoyh02OrRFkWyIWzVKL2mGH9clc+MHyNox85b
51SGfwC2eDxwQBI5hYBNCtGlaITwWDbLTO2BCQOruJVisHhdw/1oURXhS0pEEu0t8S11pEaKPg3j
sy3bKgufJLMhCW5f99nPW/3wgzKwxg42loCrhLowtjVwtG3JwXZJPzPp3hwVlh1Pk00jH3VpJrjZ
WFa6hgDHlQjCldxyHKiP0JnWEwoKRIK00KNfhZoDK7MkFhBiz69q3Y/XdFLa2c1B/rivREhBWmMs
+d7l4PAkbOJRlcU/ONf4GJzi5HYdh2d7m9gg9W4NB153TDc8j2f3pXEdShFb3369aVeLJjXbZbjN
VTavR+skGEcnp1BxZ77P+lwWgPDmNWbpqXUYS8Q7jpNb5uZsjapFl9RbeTXRcbDzCKxEFLR3odXQ
h9gOom4aAF9H0DyiMHI0/xHaDaFNP5Y0eGFVb9T/QudB9G2eEzgSZzChz7DIHuaBPFCuzkMW/py9
B+U2wXHlhpneBlej4yyqHyg3ej/TBLP6zc7fEF/yMdMw6g4c8c6LS2149kl3btmRf6r8UuDSOjbK
9Dg73eY0qRFvDQsPO6m93iRqVxm/4XflfMdPTaToWVfl5AuR3Q9NyhP7hLCmvQCxZNvz9y4iD1rh
ZP2YmViNnxJ7anzycMfPkVNiSTkXv9guEZ8bGQAh4cAKstgZ6vXoUbl28ZpYj8CIGDjvKLq6l4Vp
nH4cS184HQFyq//L2uvu8S1Kdisb3meuuxjxaTcKCjPPtDlL5RFo8SlqOcz11wqP6MzfyvZG1XY7
EVNdf11vFv6C7zwlOt1zLawY7lse+l7DPW/D4c6ZrF9ca7stbAge3fOKvB6JVyEZqVSXouHBuibA
pcRgjkL41nPyo/OCd+m4Pm2IAlOegdpjBZYu65bsBSP0AoNHhqXbq/Pwfb8XNJru106yZv6hzpP+
LVqduJW0aUXye6g+kULY11tJwO3K7p6qrVyBkA/hNP7/E442Q1kEicarDPrld5Gr7++eVGmwdHmX
Ipo8zel7f+AvvBEtlj/jrlZTNF8/B3U2G57OSqxuEXnmFV9+qYew1IrgoDAo7MiI3do+LSWdxgF9
8i5ByEcBJAoiU/DWXiSNF11OfVIZ3HvYXVgmue+y2WsUlcltiC2J9RLq6M2cJpPWmcEpKgNhXO05
/Outbzs5AMpQMF3MsPY8fNh6Cg6RZUB84Dyaja0NFs38YwCaGgYWQDky8g/ELzluAA9c96DvAtjs
PY+JlWquS6SGjm4ZDQnBjzUcF3J+LlqMP7b9irwEeUuhwW062ctrXWJxG5T9MFeP9FDHBB1FUr9j
kim4t23iq3UIWDNxeL8QLe44kF0quO3nnLJ/Isoh1o7DwpnDsbtMPAQMYct28bQRN6PzyhMJQFS4
a0DS23odXApIv76SWQj3I6e51S2Uapqvcx7UN9mYsDzDgn3vUxp/CYSlh56hht5P38XZJfUH84xv
gkSNXx1u7FiS6fcND3qw+Cpy4ZnJd8t0jjzAoSgVANzVBp7aFWyZTuL/K3cI/+IsKLlO8p38caUS
n5ud5jngo5mg3n/a82aK2ZJKIoG9qeeEXjvT7ZoWZJvhGKZ5KzKQ/yuhgzFD76qkZ2MsmrAjIk/9
wVmqJcukQV+8rCWqaQe29LgXle98TW8+9SPRlW2BnrGnH74OrJKfiQoLZFvxLZsY+bVTkGbB53IA
g1bnTJ5TQJtvk39Wy3VI55o+Jvx7y65agJeOuAt7Azk8HCASbxPOF0DJ7T5qyLgLFasJwYikyATM
3APd2b8h2cyFqq6aWpMJk649GbS0A9qynaLJ8DNh79cLP35xxYlD6d0+3azStw8980ma44gb7cs3
b+u4YrNWYhO3dXSYY97PNdcnxNvnz5R4e7UnhzUvcvP4X95h34u3KbuTvQzqbPBjoY/AfvDSV1N+
9GuJwG5ofnXQp2zSYnzjPiK7RW5LvMeKyV4vDWBkXQxd8MpObXVR/WUjJePS356luxAUfR4PvfuH
hDuNEgYpg0sLSb7On8CuAGgaZWCY8K//xQMtFiVA6ASTJe572+8PXrI+hyvMr5ZL9oMXiTeqw+Bd
8bl7nmogyaLpwRE0OCfWHhkC1qfIYbauaIz13A8NdshIkhmFtOu1gO+4mkwPyBXazqnqQsuAsTYl
ZL4+df7L/lClTXrP/cK64VG/jpekuCBoQQzb2hdEJB1EdbV3XYxhXScTBkVRBi2cZg9MwTi1wqW1
Zru5p2Ikjg6Bys+TR6FL5Ewa8fF6iVOJbA0bT4979CwhjjWpoMC1LcE1KXjGehlmritq9gRCJg5c
yL4bkgDS9H11pRRc7xZ/J1Ye1Ru8RwYNQ+MorM1ERCiBVhbm+/kQkoaThGrwL1+xS3tnLslens9O
qdVSSqCDM5cGUDjb4cqE8lE/0dQ5q2aNobEFOWvYPsCGxVaSADxynGfeTwu6UQRwlyzsOwnysKVs
4vDcAZPNmUa5zy/BRfNWdeL8a/mkLsudqvCVv1FA5sMrleC3/3CzeVbW6SDBs0zua12VUqElGjh5
7F5QdhNeNMd94Zw7yyZOwUsc1+GL3UmrSHdF9wblICYXqKzqI4pcpsYkXhZKt5wdxtIgNDhAb5aZ
BiMMdSbMPFwjniyUdG8mdVRywXq/hH82G5RTpaL/dfWNQMv12lmSv8BPMWLeRHNQlEJGsl/bQK/O
E+ZhdX/ykQFmgMjC6uyPfKxzSo8Xp5V7B4LAez1OezdTMvvB9YzGVdmZqGHfWyC/1wsnAPXd7c65
Yf5TdHCb7GHS+dryd6CCn+ztOE5227zIzcAqn5cFjdGqKSWEkKLEOof+nrmJMOY5/kCAtJ5VbEiX
nU9Dv8wuU/fjmtoZB5QHOlTC8Ktk8UwrlXBY7Fju/XufbRltZyGBK1KcQYbZAD7B+MDTMRD0GYZb
3y2Zd//PUVGs/LEcR9v6t8a6fzm8rbseYtZIkX/ILbrhP0CWAAXSB2WB0nt5Hxf+5QGSyUPuEfOe
U2fQ0cqDahlmaa43/7LhlVAQBRqxFlYMG7SoB4TFYhhByPneovm2zIezIHt5qHCfJl7UruoLFomD
Chik/vEVYK1lvlgBN3W1x/7Y3gCLm8BSC0SG2iHRh+NTyApAKMDNwSmdqTv7ArRh8QEkFnDz2v6D
SeOdy5UQ2kTCxkefBbret9bEFjdLiSAyVkN6XWP6pdLAByKueFleUFXp6wvZNQgr4xUGQ7D9iAGJ
Z5m9Rm6sLtAD5WlO7ymUVru48ADowBWHtGK4hw7CCubbpk1KZpXUs1zXNm+o5zhYtTLcVoisGxrT
/mKvC9XTeGle4W5cpTxVj9gdVccoYzDJFt7ccYW0KhoXGF4cfk5mv+VHv9BLEq1fA+iuTUyTYVSf
YznXLDxOdmn4GIK4dcUaXtN6bEbfSZDcfqxkkCWK3vPNaMr0Yo/YhmWcpWFH25Uc3rTfOY+xmBi+
flS1w5XGnj7x8SxfV5KdcAbsCR0fZxh51hpakWHca4TkCLO9uib++oEVCLHz2mqcZX+cMqI6rtFi
YOpLcIDSxXyuN+Vv1pTzfNQUDTMgvJLpHhgjtRzQZNx4gUxtH54uH8tho9JKrgmhMK9thZ7sG2lF
30ZWdpqsVC3mehNGBOaWde17doDJRLzdCPm1HrSdwAgJ50Gk/GU29uBGxtZy9+YtD7ZE/3RHPzmy
zBjZ1MOfk4rfghqNgE+3EEHgEUqAQr+FkTyduefKi1H5ep34gPtWHdZIIMKi1rVZz7g7ceuEgKCG
9MX6XYlmaQysRPHGnQfaoax5NlButR3PYvD5yFXa8oeyavxB009dQqUFQwbDHreralIs6w7/n5oz
RayMLtJ72dp7+pFdzuCD19eqgMUTfBIsf3mmMEjt7CSvsDR6EyrdBLvM8b/ZEXoBbYeUk5dl0BB8
ClLzMezmXySkiJxjSNZqfz9i8eHjII6Zg4L0zDamwU3bk+NNX2uDSQUckrY1p4ZfHZ3IYitbZDxR
pV5qi5f6NDgLXVJwYNFIwj6myXvDPPYe1zpQpj7xF7kjam870vnQrW7lYPUlvXaKVMu0MrtMmRuo
i9/5mtekF4C0jXG5VsDD7UfQLJuPWWWd/WSNB4QXXYI/a3m4xz4EeYc+5o2K6B4+2CVwRSERlEcf
Nj23f0VkMEAuXgEk9scLQAO8+Yhot1B8jzkDreWqmWS4fwKrompxNTK8r469g/6Mu/wgdawaH5Rj
KAhFJmKzxyVj0l+yo56U16vZ90/ZsND1Dsc5h1LHMo0UvTrsUkioO7YObMpj9/C3BRYgRjkqjb5o
pE8TAXBQ+tTJ2Ux2hXZgQtmMwmlOrNd1eNFkUyqngmJphr7TN/8UK9g/QgOfLyAzhlX8i75ksFRa
NPBgF0NFI0QBrT6rYWzppLQdP6s+0DSUkG3IgE4wKxNSxxuyz8wgnvrqkbsUoR6kLSPpwMmFJd8D
oQSiPioziVj6UAU5sj7fpmzdE7HdXMrTwSoQmd//IwQZE8llAKK7nSAI3ZZQkLh6DaYWHj2O9xCB
BEat0YAiDNUGGEm1etJiUedV7FesDoQ3HLzvIObLR2I+Lmh8ibYKXnWWOiMUVXxylzYU9CQt0Udm
Xrot7FG0tdrcUM1DbcV2JOjuDwnKMZ/ES0fsq6iJq3jLfJbhJcIOOcJ5ZjR4Tfx8uaam21BDUm5c
I1AFFB3xP3V2cbICR6vz1eAWmW7Jvs8FY+X7pMmbTdDuZGp8XP6qJ+wtf5Dpky7bAve2riU37S7v
qaRBSOKDDxjcGwFeT639ngATYpxbZzzqdBK9LWQcnSN8G3Vj2t3XWrwF0mF7K6walz8i2wYPUPYP
GrwJCahyiAWKnJIo0ktrSRdHf3ih4JK3YzaqWpxVGS9ECY2qAhdEY8vMoTxqfF7xKA4LpIzdubOf
GRLByjDdS3usC+ohxCCebKeYRNh3H0xd7KwFc6FG9w2mrFRKT+erKr2wV9ECE3p0+kn45hZ3WRrg
cE11QQRSjHRA5mUPV4uHkhH3T7U/+UtEEWMNsnBgqp5JBD1SYTflKmrbV8gJMG6lBqWPMZFPUaJX
UjaExTA5NtPo1wKA8dN2TgsVBn94BfX83Oj7z0WePFz7LlIAhqGk3FhrdYLlB01B5367Mukbpw9f
bSW5jetcWr+hxcGDP597PlgB6mnw64afbI394GTx/OTAxaPdYcYSQ8upXOfzSAJ3uvBwCMwXmUEy
Rn/YPuiUQFoEcfCDpeROZrA3+CHrDXA7bhPyjL6a15vyBGkpOjHUilMLlhRhjtuUABAgn9DgGH6I
r1pETwbsMPgcQAvqgwMZ7CCJ7+gyURACfdRXRAUPJtG161ztig0UpeBghPwcFKVQAtN3FtnR/TUm
IT+ZC9RMoaGWUCM12Bc5daIdSXguwGWu0NO38nInB7qUOJuawQU/qGA9gW46agIQhUAmI8CLqi4N
STgOuHtTODq3fvIlzNcc43rkRzeR/YD1JIypaldJC3/K5BBibXXvkhWYSkyhFBJ3GPEaZoqBw5mO
2VNV23OaemQ3YrzE9AqDpgPOq7wX+5BTy/AjiAAkggp8lZyIL2yoxor1Q3Ulco5AtEEjzb1qK3hI
4a4CEgGdXp+hPFBdTcCVjAdCU93y/2Me8KWvqOwStaoFU+NYlMYqRuX3j/YJ7G/iMhAEa1PrqxJ7
wE7cR6pbaghpuWdOoEKxP1V27KcsMV4qOX1AU2HNuiGzcqCZBprDUGu/IYKl9hrnmEI9TaRYmQoL
Vqxi0vfTtnqA5yw/Gmno0d824x7ambMtpOJ1IAAJa/TMsT9yYCBxUk3DwEIfPa1qW56q7QF36typ
yME3Y2IEGOWHHeppzMsLyfUH4rKPvMXRWAz5iwVJIK8U0P1RE3cpviPVeus5n72ddlyPrnd4bXPJ
5Ad+VNC9uJxhdJ1tCV+1REH6U8iUUa0XX96cLemaQlvDSW50SeNBbtwy1Ot0n9ImhXmWvWab99wI
Tnn4zTOPlvzF+eL4YzKljEgKjPCJy9OK8mHVjEIUdROF8vKk7yf8fuEvILH7WY69rIknkL3wy3NF
/4ZgjCbhO9HUXL8IxZOjiF1mUGIZF8bJxenC/3ksPBI/cAYJ2cW4Cr1JHvters6b6sfHiX82FkS3
lqCQNN8RIEMJw27nA7xzxTcliG7nvxNKfiFnG9DjdszMSAtx3CUKxZIVFVhOOeY5OSgTAYkzICrH
gV0o33HrJ3xoKrY9pnVjRwRtJHop65Lo+cu5vtE6RIH13698zfzREpL4t/yipDzDbjU7Ap5/xdH1
kvo3Gv38hkqUuQQg67OVA2AZ09HzQOUezVyqi1CnP3YSs/rTDnGaaYokm2VF2GyflgAgit8fI5hO
+h23TH4gR6Xml+zZzNRS0oBO4kfEDJkyS6xJj3cvk9w8wClevHLgJpT/6Sj6n/D9N8yZHblhjkeH
Eat0Nst/RH7zfar8a6hekoDl2qVlh8ASbRFgkyHnvyuzXXLaXjleflDObHyHccQ/HKoFp41zWN3g
IRyF6uCaZIC5fDplyW+kqa0iJtUCILOMLo2TzYcGK89CQOegIGO9IsiTeHAXCZwlN9Rs80j+EmjB
m0aBixusOWhSA9hVO5ASpasucEZGIVvBGbEUhy5cpBiMS+AP979YxoaoXubhvxmSiwZAUbqeKn/+
7YxuG8sUHmuvNz2XmbfrWY8aC2RNaE+mO91yOTnI6VYFBmszF3fL8BetBXHJM/GzX8doZdwTWRQE
DMfKT+oEhDdmgFbvrJDf5aG4l355BCx+aEeXaqLwj8uvpbn/1dpRiZ9pVn/A3mWZrr8kXpl5pD4K
Ege75bIBPBvSJg9y8EKiLyYVMJWfL4PMySZ3CrDG5r4aEDP9T0p7DfRGidcSRwM2RNrRf3jrX1Rp
17o+oxAtbYDV0DIt49S4L6dOKAe32oo7vHWqqDpVyk+35qCjAcRdy+ddcGJWV26oCp3LWX/b6/YA
SfJAJPxZUTUsBaKsENEiX8JbIa4XhldCNpUIvUGl6kkOk+i9Y6aCgVzmDEP3azGJHR9VqmOZa+3t
489itv24IoDddKxWDVHNVPtmU1EJVpsbp1B94qdXr093cb/n6tLrq2VuasY1bPbL9efm7hh70KCF
4+M2270jSe04ddAebVTqTfHlwVFw3av2yuMVdA4apLLcAQmijNKN+TlMN2Ast5ApRo18ynodNjr1
5Xi+7YrvwTs14OV6erAczgqX7Kq3pOQc8IRZPkJtXDuFR3yQoK+GlG+5KYPIdk/Rd1S7T/C72Eu/
cOlc9qODR3N2MzH5F8/ZpeY0k5I9PjaVtcucafrrRanORpSQuV7UJDHIPtc7C1gGRDgg9vRPDW1u
SZyZ+tSbS+dWfSodotVMwVpONo/VgLu1wkI0iknLByfeF7fH84JPZpu69jPEMb10glY0Ayp4lvOL
UXeVt4eBlnUI4PwnQzKOHNzkS6g1+YMHxr464JbKm4B6jpLPGFCeXfm9NF5ToyZhPhqsXhoLTaUk
/yPd9RmoEjP3MKvHhBevwwd5MRBJYu22bXCMNL/GeOzddUtkjNUy7IfeReKTHlf1ogg6G/rtER6N
E9MArl7Wyq+Xk3gofp45wB64FHYSBFtc7tPCLxyqDod8XAbQk2BmwIbpuw3Ezk4IpppGZKtgw8t7
IRnGOnA/M0+P2b+G8O5V8ALZy/Xkiuvwi7bnQ/kdi2dLz+9h92HnZEfqfaZKekJoeg+emoUa48AS
6Ym5iTsLnXUS/Aq/2w6ZINKLHA6SDv/qJzahSZ70P6D9NST3Ah12gE4gDDDxipd1Vfvy7hqJF7s3
BcpDkuqOjXvjfgWr4+SPZXerRILfVxiXFhaDhjw/6j6WllrSCiT9RtTLp9fRC0F7it8FHCpoJpuV
dIkhhkD/GHiUJNkzNC+RnsnP1ieT2pZ8oDr2IAH1pGcxPibAwEVxt7VHXqlDP5SvBee5KsM7gE9n
IwOuVFBHXZdXoDhT6mTpMTOWPRdvNF8SJVNoKs7SFD1lIbV3e9h46w54LQ0fQxQixbKQAPwX9MUF
aY0Z41KeFRXbWQfGlGAYNyyuT2241+bk3CRq8JwhGFZJz0vM5dfS618Y23BAthn4xYLD4UXbXm81
gfOlozZ3JuFvglmJvnHrojunozbpeQTV1TAiX26YXcIr7Z6SnnIN0lNoaLqBF9iJhA86H4bNKr0O
eZHlif/Mt1zrkjd37D/ZtgyHtfqHyEPL7bdnKjAXT5bGS1Kh8Cf7epvyrBgGXopXA82xvv8Chpmz
nvagjEP2FULvcs9fxzXRs9kC3Jo3+hOFo8vDFKLOTB5vC3+1PTamqOiyAGsDdvV9KLuBlkJ5TbBJ
T/YWULeo9bQtW2VGuhzZTGhTUbhaV4v4KOGALjEJHALq6P/mJa/JSgNbwNvprOpOPjuIzVNy1Q5f
y7EN3MJDULQYEUDIe5UD+k+lxFrKqDxD5D/W77oC3folCgOR956nX32Dcd8Y4gs+TLSXCp36sppg
cThRrFuEMSObx2lMasCBKqB0s0POS+Z44yxVbBxCclarcsr3sBOvX4KOu3rvrPpMUJHeGxog451C
ejQsklDOlwwFgXAxjh1xFZ65BE9ISDiV/6uFnsofXAlxThjotnqQFwDEv/Y5DIu5nPmtLVRhZGxz
3od9W0MvYmwtwVXt5f0Lt8fO7C+EuM0u7XYgdr/Yej88GGKdGe99/KiB9V7cW4BjWYkI2qff9v+s
N+GnVLHSy9bFlIyBK/YnPScD+BJHZTbsEpxPa3LbYvTMfm6JnmcHGsDGb2Ea0sfASRXch+lZleQT
Zrrf9QszrSFeXHRepLKqgNmlGQB0DkJ6Xc/zJaSsdfaib9Du/LcEgoZP8rbohX0l2Wdg3xw1m5rt
DhkJ3ehW4DpHfalknRsacjDtO+ZhELsg2hZ0jbSnzRBcRtfZZFw15sGmb75vwDeeifuYCveVVnY8
aTe8InaACJAvPB9+YC5Cy9RpX9nUSy1oKaziwrpMaluxCGUI7omRWja5XBu8c59ghPcDwHzdxVw8
EWTFYssaaT8ZlhGDI/JcFF9RDBnP2Vdjf1RQ0uIujYru9ywC4xI3q0QJ6t9N/m5HDbj/d8L7nNCb
6BGwRvSitT3gBnfLm0I9po+lLjVZUEva0FJqJ59DEdbnTNajFbjul7xlPUXs0uXbp2srwMlwwyjp
gZPh/1Gfy35+3pRkS7TTyTc8GfluVzCEJXqUP26DpV5A/O614Q9Z0CkCzQjDTahN5/oJZhF9gGXq
Ic/dXWo4eozcZWywVBz91mVj4VXOuDvMYeFQODQAhLulsKMPK96DDbK4JHcfSxH59KbqiArbeSGr
aF4fq8RLFelyszFus0TmxsypZEPkfkasLhLvNPxi9fg8Rit3hFntp614Z2x/DdVauqJsRWiK1UKR
Bew5v59d6Z+eDNQFLZD5tLazFPrtKY0dCMW7x6VBaSvS1rjvbZCR1k26rbaHdbjBfkvQshbpOvdH
Fcm6wn8A0sVUcuCqyjJ/1EW0KtSTCEq14BACBY4d9hrplMCk56X5MaxkM3twXaOx8PsLuek0lmr5
5qk2A/si2rA/g0jvC+AODG0WWlY0SiIXsYjZkpXeVf6QN05iXiQ9e62JaZ059oGJGa/a4++U/6RD
i0rtJuZDDB23BImH/H6Wk1TF22rJ7jN9nYXJjRXcPPL5LZYAx1H+BUJwajIY5oh/PNAnVZRqmkyC
gvIO050cTC7u0hEPYtGzPWfrZz/IHE+VRS3rgwx8MK+QdJ8fWy7HaK8dDSTQ9zB51tE+chHqG8FG
+htv11bT2anyBBKd4fBbPfZjIDlAGdP68pLoY3IGVphrv5xst3XnHxcG7AmP785ju7SPwx3d3Ydx
SPHxHpCcADZxUeO/K/rBOXirvtlJKTnKOfzH9e8km/FjyVPMLEuyBmhklU3PsFWEm97Vc7ZpCN8d
zLc1dOIRkNqOYnV0wpdDF6lJyPcin7CZmVPg6R4sQm6CZdSoO1mrjxzbfgmfdkMCTv7Qq3ljgoqx
q1alysCuga0E8whh9AD2Yr5hjk4ZDwMPe2BGj22iT0PmIoOL6s0v0DmjQO+IOuTpDXX2BPMzS7jW
gP2J/UXtQSh3KmP6KbuC3yiuxQPvhdDMVh+yilyXEots6ZITtNnXBJe710FHA1Z74lu4hTiMOY9c
7WflCZdQ/YDaWvN7/NFd+BRKXeAAIjUnNdAKGoPUdkhNZho565lwswIhNjbczo/YQ9MsgvOVNiPA
uc2DjF6jKPrnBBvILPtp3L3JxeW0VAqPNgvdTljMY3+odgWk4SFoUeJJLxqKwtdxQPEheHk/BqNE
dRjgJ/tFWEn2+M/9iG6U1icHsqJjloO7V+KvKoNZrR2TpJIz23UEmNN+J1ebYJaX3vw580RN4sMg
qah98RCA/NmgFIP6blG1lI1qeXd249/rcWFSaw9yJ3mtTIq5jXtrLtGsvDibnbi/P8/tvRTSwgbn
CT6iJ6ujz6ht8ApaJXbsvY4k+XNtdbLK+sni2q8L++6okgO1Dty22IUuOEXhx/JKVaaq/bGgsFNw
Ed7GIi5LDBJM6+UYBKUmYrR4sVY1E2C8oyJ1Zq984yAiE7g/1QdBKV/KhdaWccunxPHMsxfBacsd
nHNFf0MPBP464g6Ejx2sGjfXBDkM0D/SAxyftx3VJUjIKi0nvTE8xwiRpkOIODk9zJ9gTVr0mlhu
+/2ja9sJlZsfcThOTdisDno9YcxwNQtCW2ujTZT3bN7u8un9TPswX+lGZxIZSPR2hIq/eGsP8leH
ntGmOYEGGfIAOkkfG9Fh8BoOE5dDxB/ixPWQP2HuNEYW/5yHT00JxRZgkJ2E9cuU+Nb+KJgnLS4F
ykAYzjWENju0OZd/tM0dHuhcx0GSpcr+zBPku6vsjuMV3RV+/TtO7NcgYIS83m+l1TLqzLQz6fIE
K2e6M+WTI+Xc4xuaMnMvT6Y7Vzil3C/TRD0UVt/90wTVzvmuSRwQ6D1yovs3dxcUlDoMmJda3dHn
F9IO9G8KV6bC26/iYfJko/MFHJHbPJM6xz55pBXUNYl5yAbplnevlK0oWeBIrqmYP0vldho/itTo
l2nPNG+Ll1gdtO9PbOrfVderD7heOPIYvSjkyHutpnZHHnR61InBGckLgx8C5b9Nn5RO/Advgkcu
Zl4JZS2shcSafI+zXekZ92fcGaNOYzcNs9biBUQwMl9lYDm7cYV2uf3nbAxld4FM6frfF6n9c4Nl
Wg74nIOgqv3LmJGD37Hvn8aHw7sZWLcM8HA6HLjsvRDI+QbsynZGSa/PzmMkSPDhsazyn/Lbxr4E
b3lRANWUO+95PoYj8TzY807ekbZ+btlE/r2Ks9IwyzYSj6JUZvGJ7D7UwKt/l+OX305pWa9fPFTd
/N0Os7FU+sXirFwPeSt85WX3Y7R1NFn+uORFBy9OZmOhUIZGENV0N1h30IiadkdFqYc1iflFfaOX
zNW8PYdWrrX79Bnb0oLOyyR6qHp+c56RzzsFAcSCzV97Mw1eKuPPGPpTJzp0BP/RA6AKi72z39RF
Hi38gYm6FElDS98z7pbbycdzglJCk8bz1AnoxSA2wgh7u7cdFHD8q+5vNkTS6lR9l9qU3FirZAMg
X19FcakNue0FeJbKn8ehyAxKCdjFF9OQBIo73wNYdA1rOKYum4x+e3L3up4MejsMtcWLnYOEkNMr
TpIyZ6un0SEXrWtzrFpwYNxURBBRWAcP/ycRWE4ebmpwquyprZgrZ3J9ofzfV7BNn6E/iuyjo6bP
awL+scLPg5oXrePz0cN/UNxL17zKlIVKcfNoN72Tx1GYgHsix2ui2FLIeBYa5Xf9PRvJJhSWSwB5
7fZeoVgSab1Zfcbq+ggxKl9eREvP1Je4weesBk/Gn00DfWrQzMM/1YRv/hQkyzUogYBh5jv0J93K
XGC/+pTPAEMGC/BsbeqByp2a5hDW81IlRvkD2+Rt+WrKRTvNIItUnF4BSRkWvYYA4u9i/GyNfQ1a
qRY2UDTwKzsoPZzOWwVMUar/aKlhXWjvFLAuH0Ljokr5DFCG4NIr+FK4XKDglhrI9WxIspWGDn+S
nliH/q53dIMmKNnNEGi7rIkI5BJUI+ZatlbX/5qcAVlTaWHSiGDHUfWSl9PcbnLpeBGkarY2oxhD
OTlsREQa88Z/7QXV5se3Tltief/0afZuFVZAWPmyEsa3LAKVJDhZXENvbUwJwkNxquJ4YVXPD4vS
/HNaiPbLcQJYE6i+FsLmuPXJi5LowkGkvvIbCCVbpPaTNnn1k98rA3toNV8QP3a4V2Atab73hyRp
AP1kCYMa9/PbBdtfCp5U5usHTFxNVkKvJFT8bX+SV4BphtxzCqjditgvEP1dfGixOTBoDEEvlEr/
4JmLlhsOtjNGFYorNX3dKTn2DlKa2flSssnlBo3GZHhhDNyx8S8B1fITMMN575sDBNM76d7zJl/q
opfoZMDMk8nMzzD1QUAOpfrfWA/NfgyZAFikUkOcMoT10+NEfbbu1+usyTL75YYnUGV+PjU5UcA3
nDVSAtOxgyeDM8fZkjIv7rpqaR9hfF3GfbCSlyhFzJCp7EmJcJ5PBYR54vXh1rcaIXeeWfC8wJFt
seKuNAyFqI7SpXx6agMQlpE+SnUKrrzkjd5MoeXjCBZEKjIz9NJK+mqehlxbn9h9AXzl68RCiQdN
ml36kd20eXENXYh6WfaAAtxciclLezmitnGsjDT3kzgLFl8mXF8kIzJch98tIPbHbX49lE7DzF8c
q8SlUj/zwPZ+YaOO3c3bTcUCSJt3tN967bWo2Jcj91IO3lvRJ8oSr9OvBBpCB6jhmrb+ptqbS5ZS
6zHsbFvJQn5YHXWuu66jFWqZZOIusuRbbGZNqJx09jxwIVlRcbhgnXe6LDWYim0kEAIj3lq8Dfn5
uKzRBC5uodVxbts2fKglXeZTwJqP532/V+7ekvyNZo65WRiUoy+2rpyxtsLrW/kJuC3vgOhhcNef
zApjVH4lUXuqBfWWFTRdUj+5NrxaQnWk2lVn0ffkvzLWrYKnZALwcVVz5b/34HQDRNGrD+lgXaqX
SCP9Iyc3H1koydeN5qj2mPwa4R1I2q6z6iziGk/c1cHRnZi4vABdR7UWUugjMQ2SIX9ACPKDrDCl
jRE9L8sFseNTb7mJN7cMfl3uEEZDPgF36bdcFVnx5+nBB/MjnOc4n8mKzbCxndaYMaZ8XLD6cDpu
DXagQj7BWrbNBYL+EOHOiLT9YfbZ5hO2yvBcK8CxYTsT9cFtgEF2Oq8fBUslqqDXL0LXSsRFTgIG
K2HWG/H3FX7ClwQeGEz1KrPOHUJS4gfs42w3/Otc51HX5758C2QlCAAL1eSa7RiQc8OfNGeJt8UB
dxPkw49ewAY3KMuZkkIUznuhdFt7LzTUpjsxdJio7vBzB5DMl+LDBYPdIeVzX/CxcH2+rV+f/ZjR
cV1Wk61KmWpqu8RsSX7aP+XvgY/XvWf+01LfeeFhBkMVSDZP69aQqNRVqah78lWFgktW+bCgIiha
EF8uUT5KjnvymSK+3s3pZc1oTGILzPFv15vkCUZCGoZ/a9nfLGAx8eEO9S59aTuA9IClvGwfR8Z7
4kLp0L4+MazS9v5u+4++GdiU/rHvM72RBuaW1oOurCCB0hdBrheva6tRA9XitgaxCWP9PXZH5Qq0
VeDJkYnFucOpyyRUFMuxL+Kj6+YdtjDcOpyYduUEiN5O6Rx++2atOcvtokCOpLC+2hzDLsGCXHF0
JDJEOWSxw7oGXhygNrrWIQDOp7cAN7XKzV8MdpnI7i+7wfsvBMb0mQ/bID824hnwHU+xxzcy/j/t
/X/oK3lQ/2YQsaQYBnmQ7IfGizQGKsfjOwXuOIiYdxWvJPwFAMT1VLnHqPKbkz2fdZN48iD7/xJk
+iS+NDOl4uZ13fk6VCfQyroKsJhdAYANAlpwqtdgHcycHIoAmWQojhwD+XXk4C1QrvKzTQUVxZEq
2G8Hx3VhGl2Mp8y6NzUVdsEhmWcI2MX5ACZyI33CVskOf/NTZSGesebpS7c5zh3put7m0D/XNK3H
nD2OF3ydbp50YIt8Op9L0vl+iM2ST16Abt6dRoB3ARPpIgyjLfKkxzXBumtuE+k2RiKmetZchMDH
SmK9vRaSRcyQgUqgo6czWCe4i9CQDMP0NgJflYocPCsJ+D7+NyXZr7+Q2s5TWXiews/3h0EUtQ0a
MUpKyKypenkL1c1vxsjIH/BTc+rfLA0oo5vcGPfbH5YwJmJPNBbuta8cYsib/dVX7BeMlCTvflFs
fNJ2lFQTIkf0NEwzmDnN4QGPYkAr+J67F9MfAf8YphARP6PBTnDfmgWJMGHn/4JZ+x05qfWkN0rA
s92W65UqiRuVV1MkbBl4vO1iyW1ewbY8o2Wuumzwob7pfamBDbqniMTFp7nSySsbcBoB1dF24cqQ
J1Qp+eo3Cl7oK3plMp4oVG0kYoGpnZiATr8p/0WCwxQmup7LXCr6iIq+pONcH8uGw5kCl2uUZ76d
tHBT2to5sAIZjaqkIdGtZ5ck7QkblF62hBY2HbkOBZW5LhKzRWwjvSWiVOv5RjxISM5hPPg+jcS4
5/WlYA1b5YrGAYRKl5/l9jrVsAHSw/KEX54xqYYBG1eFbPIzEqF0f1x32u0mvxOVx4HCRjsVAoK7
2X4suULeB1H8CvyFYwlftLXPlR3UikuM70VMOMABdmSIDZcweJhlhvWrMqVdGfAqM24hgfAOZFLu
9j0GiSXN0OvojZwVJ8b70sONkTZI4P3VXPx9rnCc5btVBdBAA16SvxD0ZDJyrNbiigaPfzI3oHA0
w4/gWYk1jL5cWLVLKqAhX/oOySxzpYQtgIJZnpVv9D0+kk0maXVpitdZnuTuv3+kmox4mWqWJzlK
HJSP/8XXZA+lYQsJVlwiO1aTSVg0lIu332foi0+bNATHXtkPBxHoTJHwhW+iKJPVYL1fJOb2m70N
cmlIajHmz+gmqXyeyGoXa2Q3rzMZsrx97im+rnTKMDid6lWdbmrkaj26QaMpF4AblwZxZiT2/pFx
uMllE7TjzB/GWUYIzA+rgdPW/OPCt4QnllJ5e46p3SDWN7zAc/tVgIruvrIN2EeJFReH831RLqsF
h7rdABHXnwud55dKnRTrxgvXntWqmPOAqQJ2hGOc/Jevs9JGirLD6e0uazVum8P76+UhIFQPbqZw
j63RYW+y3cL4J7LbeG2dibFeEz6OJcNHc5d2W2eFFM02T4nosGNs3UeVEmG4zdCdKx8JotxjjIkE
6m2vgECyqqgYoIrl11FIPc75n8DetH2th1kGXzG/9yBEfrWlvrhbGwAHHUE61Uf0mgs0RQEPMayU
9KtLgz7V6xTUSFn3bmOpc5a5sa73RuKw3YzyTQyrr9NqNPdjsZgXRPxuD/YbWQyHc3AlQcIg9CgL
MIPsEHARFCDCqH1oPtmbQan+7ePz1KUNuD9hElqfLvK7GMS7LmGGzcOItjo5EOyTNdb3S6H19zzy
zgmgG2JufMkzHauLJ0hgYevDalkK0LQEGA/gjtia7buoJ2TsSYS27t8ueVLYNb0/tr+AmuYhplFq
6EaEZduD6d/343HpjmWfhR+6SqsEAfj/u26B5QNhiHVEOtnJ4nH1i44pv2gDfg7RNJ9+7tUUmqlk
R6Y5PsyISJIiFcmdJzUK9tevtBbk7MV6YfhOXTrEog+0tbDlj7vUMSzKPT63I+nFgFX7meL84uvK
j5+DujiFN2CR8CvVGlntXtX+5SAfiXiK0gwOtTErAUj05Ao5+x9jqyNb65LcqnlVbKzH9wUOEXaQ
Sx3A4sTjTmvAMy57PDoSLbPmkFzmSr6rB/ufou01iv+1KF1ZVKrpaLcMsechM52cC/HvkMWDiXTt
HQj3ohdnAWJwqOR7ykiGE4sNSYEcTsvAjs+ARoPhND1xPoMvV5ArAJxXT6FHHpeFHKXRzvRzdlUb
PZd28PjCUB3Q0rkNK593oRcKFG1i9K/YmYeg5TZ2vwH0JieZt8FQBuCr91s8aMzVXC1HIlfcdmHx
Q9aha/pvj6cf84N6hMBdOSrk0DBaoRP3pYlp91cWnuS+NLeYlpL362uUUVkcEWZ+I/OhSoWKjZIV
hJjj8qqsthLtUnZV9y+c6jCM1d2hIYhoV/gbA0Yo5cbHNjg1cXRknzRa3ItUEpY5WfDFecurSs07
tamqABFmsJmGAeEDti2AooFOKHnktNiC3IGKRrh/Q+eflBJ65SlL3M1BERhejMPvLzE79XwwtcyL
u5o3fAbymTtOtZWaRvFQopEZS372MrK5+mIDVJ84l8idQ+quLcEoPKOcRKxnXvbE6HNaSZb2bl6a
Okxi99Wfd3MB9z42yoLzTG4aG64kHOhyhCXt047cp7HvPIavRGry4IREoHA61H3x3rWgCXwfmp/f
fU5IwQsBCMCoX1y8tzQ06YhggvgQct4ho0rexa2Fu8D2UvaJRHfJJj9WMP76tjN4nVFH0A6awcWq
7Q6gSjH7lBBe99zg/pFuR3CPmtGjcrd0EAPfKnDOUWKy9s5bT7+s5WAUJPuZ3lxGAqbIu9Nbqd8h
OY2eRlcQJWjkXdaB3BnUeJGZ6GzLup9UErr7/Mpb3HQgvvLWO1Uokl9OIE+MzSQIKP8RtvN4SZ3g
QIeGnTlaba+czh43PqD3F6WLjr9mRijcLRMvAGZRN5xaxze3opp3H0gp4LJbb+otBVXGgEfNgBkZ
v0YNWSpcTX5MtrNjOEgQcVIdLQnxc2omXd5VC34AkUX0rZ4nWEu0pL4pvLRlyUKXW7tf3iZkmGX/
2q69S1J2fZnrmJEuqp86lWhj3epB6Q03D1X54DHIc1Sn7Ugm2C1b+V9ji9du+VMQuPZItNj55jA8
Qo0xxGjSpW95VoqTt+VcDlbzdxcdEohXraBhuTPbXnG+v1LYFyGvLdBYqxJs/2pcCjjLi6nc1GuE
eDmkhq8VIWmQLNe6jQ3zCMh5Xp6+vOlX0WzfU32x2V6eoTbo2GL5B4Z+fZCNUNRISJr5lODbdLbX
eVq+eeSPgOnOEFOc1FkZcv6nfaK7SYVv5UdC+ofSb2X6VjzvqFaoH2BVSu3/ZdDJqofNHa12ImHe
dzjzn236oTuv/X1k/97FZvqr8c3A7HiDqFtZD9At6Ag1X3jW00lNqUghumjoUkx45RPpdKFl8J+U
+6CRyWgeO7EPDfrTz3QLXHcOv9Cdo55vsZeMhID4+JpWorhvw3cS9W4fBu0NqWlj5iUxl4+mxSy/
0vl3Vx+8ONmLLZMy08UPa19Z8CR0gyWnVVKvSsEY8f2SNl8la5tD7py3VwY6NVWMu0ww0wAz40Cl
vlpzLZXcuUqIlZ/N7hi0KFpQq0JX2e9xQQKByP88nhvbADhj274xBN9C/1v6NI/ZCfa0QXL12i5F
Rlm4qdgUFLUIVhYuE1DPxo9/YeNj85u9S7H9K6IQZeuYPjPXgJwkZsOfGwx+UD63k+VkhdzxU2Os
IELxMe/jxCl091R14jsEVJZ6tOaYOCjPJpGpOrTfeQOmA21qHHQMseu+nVkwizlu8/fTSEbjsy/z
Sb8wod54kiXdFysFk8z6QIkXHQokhiOxP1+ndBzR4vKjWRXEPa59WYNK57Xt7ZLfSe9T5MMlMdeN
zRBAmWvBaI+KDXQ2qwFvqG4EZzCnOELWxWkUrwWs3QsgS6RO0IZeeczo45OoW80VJZzLwko2t9wk
e1hrgtx8Fw5Jz0MNpZS95OO1c2s8Nb/EgTyFNd6Utwi89NU9N066podo1jdoPdR4QLAS11Ys3JDY
Btlr/2ATsYmnPRu47YwZCezZQ/9SEikwxYsgO2ZCpv56AibUlemK6qIdjo6jo9VezXEzv/1K5TLt
4As3vKpBTLbmFYmsL+CctHXZAvGDOmY0KkPTgY4DYOwnNxr6gfb7x7SrIFEW//Qxr6kV59a5NKez
NW++bWRCWjlKOAsLFzOPlLSY04w5PeqO88FhsPTAM7B//iLmRjmYJxTtVcEXQ3G4Fr0c5SiCQZM6
Z3PV33WsxoOsVyUT7rhLe7g9FGuy30hnsAa/DST63vQQ/N0XQKA1B4s1PJQNqLXYtmdacLbe7gs2
3jU9Q5Bdfp7vS74wW+c5/UIw7f0gPtg48UlbjiNAV2BDvcrawmZtlF9g/jeUElAkKM+EaBMtQHsy
ZzRbENX+u7G3tuL1W7IofuAPcfXi0hmyS8bKC6BqdCMWw0EpCmUqOBndhIKuaiHKqivHvnjNvLx+
+LWnB1zDW/SsQxRrLSDzqNwpU6SKnygXCUzG8cfMzXNdKWk+u66tvZzkwxnc5GLFaxlEKkNxzD7F
rGrDZbDaL7OPC8RTXvc88dRIFNpaHIY36hU9Fq14dOLQUFIOxTWeKCZ1ldj5LGoCUXFdVmjPwWxB
Pfn9+BX5YO1AvDLe6i4tE7qNoyHolTAkmYjZ2R9qJZ5m34UopFd3HbbU+CIytj68cT2Ry34MuWXE
ksetAkJyLXcFpj6p56o1eufFE975fZ/6av4Mn42KQLGJ6NLyobatoTBzgaPj/qoqZCrULjAMuX3q
OjifpmTT3kzAHI10TJ/FoVjjqb/YfcQ8VyGXyvjSNi32R02/4J7osf7BNGUc4+HFeHK/VwNeLIPM
/bqXkoOr3JtZLAm4ML/HG1HMaLCOO0viKKyFFPDNyxoXuM33IZAHq0BlYX3kU1Te2A6PeiDKVNzk
lQNlqgmiYOs5+X7wZG/4bevP2n0uD4eDn4/dsOdB+KQ5tmLsrxI8uELG3I8B0nwsc2HfnxjpWo+K
/uSvFmJiqTrKJ/KViilXoZMYkaMRB3Os/7HIzaLr5+AfrH0U1vIMMTBEYkYlvV76tn99FM4sQgV4
FPxx5P2ZzKd+C+2tP/EJq+ETQEvWmnA6/TCqH4ndBNt+sN/6BQNHn8SsjOevUCRaOtFN0ucDj99t
FoinYUIgP5TtwuZGo8LeOXjU0HJXun1yQcu5Z/O11AIbZ/kiI+pAYkpZgZ8SduvQfa1/nT3bzEra
jyTelmhcdaHNdSXuiM8BEHdWXXGojtSiE877Wnn5AFpiCVT51fF7Jj5x7RKAfuQZL41CO7ERG/i1
OY0QAg0N7CSVVsyNbM6IoM85sjOKLYlb0a8vZRTI2f23pQDQvTxa4zVJcdiIJQE5Oa7CIiyuQETu
gvObnEkNxUx0OD6jrwEBzp9Xkh987+zPfZyJUXd+9SqJdbHVQmnNNsTrfXE5pmSOFk3VcvFNTn3V
iTM8/sXmv3WSI5rt/RoA1V1lQa90S5yClPD9aY7U37JwbBmcjY2mEsKtJekDPo8kY7pNWMapp7jc
BhiJkZENKRfiK9ewE9ZHYg6/nUuWGY/OtzfPhmscvDdWHKfWhn+/53/kfz3UxvWh4kfMW3Suapfl
PG9QmEGcL7QrU9HalMqFT5Ff/p4cMPCmvTwKRtXTcsGaFT1o5j02eS1T+aKD9koDeNrWM4JGh9Dc
ToL7cfkHTGtv6FSG9RPVBKBhUEmlxhIX+3hIYxgkl4bG34ChLdji2GDOmIjpLKJWPh0jCUyVwwHS
w1Ke9Qb28Ochsf0J1KN7Bq7YbtRMk67H4IM9yWP9BwaGjRPxoTRZ44YwdP/YhCtY9KoRzPEnDiBH
wZbG4FpQMCzzcN/8Q+mNEKi2bnRkun8dDJ+Uoqm0fPpanPjlU/zXNzA4frCoctoPhnpjnQyE3ICk
1p2svbUJ9XVp31X7E2lJMfGpWTl1PE6XRTDHi1UqCSZRCUGVLnUbC5wDTw5gslLP2wb2YUVvu5wV
kFaDLve+xEe9QR+G94kVSR5wRURkQA2Q7NOeTJyfbfVxldGCsNWpbGQiyOsLR6M7/VWW9ZrDvw++
2nMwULDr5zoEm/UDXR41GE0s76hxekmngOlzkgPgth8Hr0WuH8n0gbu7yj4aoIKwOY/ZLlEWP8UQ
F6kWdHjO1vLTw7Y1hHpb9f33mqKzi7bK3/948pJUYBV2galNE+4RGpTzNS8KRuiGi2AunlPPF23/
cmMGXEMKTjhwIT7mQpDozzqfpwwZvTiONN+Hcua/V4A62iz+EDyf2soWeEhYyA3UoxSAIi7sfxYt
MwQPaDu8Lb0fthqBFp8mm5eijsswhSYYWJJFW7bY6NRggrwNptmE/oh2goWhQb9rBtGrK8GHu6iI
3q0Y0Of++LGRIe8g5jMGM80/PtLxAFfxBcv7cbLc2Go5Q+zGYyIid5KWLpTcDZwaH1V3XuW+PDiz
uIUKN711NOqLdwjn2HDtNB1/a31IHXO6OdyuYrp7NJALxNjEsL5Uc/tKZ/LvAFVb2L4qjpi2patt
ZIaO0DcQQuNYeFSOr5v70HXE4LXUdVuSW5VjHa9yU/jD39oj0o1zyflntVFC8di87zGWC9YJRs3u
WqwA9VneZhLAa9ES2nkDBkNRC+I2YA8u8YOw/NrW3t6sjkvZ2LF8V7N+RDtsIKlUw6692TF1Ldwk
7lTn+4gFhp6JV2O3nmd1+a9yhLRg6xUhu5Y2zyIHYsp1SBZ17Nbh9ZRh8W6lO3ULDhFVSUO1UH/n
E+YIdWPjWoBKboZzsHGRsl57/IoxER8rp4J8DevZn/139DZw72Pp3XkZ6nYBcMnmgZLzqCirkv7b
kkFhjWB+nF1VOdalSXtxCX2QoLJG+EdbBWeY4W2IsgCOmxxY2cyhGQxGsIOX1YudrGuWNrFsuM3U
AcwDY44x5y2/5CQDllYdqWJfUhD54T7Zck9eChGlzbhijbOWfMapRsZLFwQ0H+CsDTnyjxusOY2y
Liok07q/6OmDnERPqn6exT5GuMlN5xi5tZN/oZfMHldjNTONOk377ED1T17SZqdsc7pXSB6q3kLX
P+Hj0e24aQgORg4jB1hytCiZQOY1IsMiKFGAezU1BXL01uQVYcON3jWv70Vr9bEltbfF8DmiZqmq
bFXS07bkGnz3yfaB2Ji30LjPZzEMhIg1EKwhv5r728c/CTQa4jvChqQdKM0DDZQ7BOHOGGgwM23G
YybUjtsTgKDkMdMoz0oNFiC5ISc1HxMbe2YzU5OkiAbbP3cR41U2J6DDgXTmTVXGNE/FTLPlKn4w
YgDuSQCukAf3WqmtqiRmAtb84OOvhXQYwF+Zein0cKhqZTj0KAAd+2vNS1uEP6ySn1NJiKeovJgF
iHqUbxM+j6MkSHBWLeTHsYqFcOKrwOg32Q4LLtloPCIQzVw6LwIPya3ZSlTLzvzT/8Rh37Z9xVIy
A4QPqoKU08wbJbLmS63ZOqWA987YEO8YhamyDZHm6MrWoF+Ac150RidObdXZZJQiQvOdvYUNkAMx
QhWDCkXRuxreRjp8zXJlowJwa5RvhCXuAgKzFsF5W7n745aZ6N8cfOFmXOiZcMN2LWdjiPHQchsH
WebsNovr5Ivz8DagxAaa8sp9SvXZyDpJlH4V9MPqF4J1nAcf91yq13KU2EDxCFHPk1mmgVwMhzJ0
MOdFU09jHX5MqjNekhBXVNkKt3NwhTveWBd+1i0oMGAiypQ3iyXzbpG2kcOVa/01gnaSafZno8tI
b61aOPkQ69PIks2iFshZvvaGWQpqs8pcSDX6rorYvpJQxQC5cnEU+P/nyOhtt+nBn0GZe7t1/xvJ
pmzJXlFN1JhGIjxUW3PmcmdtjoyRu4PIX4KcFBf9P232l7JVIB5hkt8In1q6ppx+M2CjuNyvCX8D
H+yMbkQ9jxBrPKUTK8yU/hawqy60tl7YQ3wzbWFBni29WX1ec9l84/t2JeCyFZGssoBaElxlZWf3
8l4egJ3aiXFwtnRnq2qT88HWxLUtP6Ia0bekXejYmvElB/0OscozRMiFXsooC3qpvSLaIMBSsFfA
+LmWA6XkWPnbDvMZ2/ZpFzYwahBDcsHH88Micm1XKMq7e4ADTlKCmmxuXBize75+/qzjk3mi/A/4
hL8yZmGDnHGA1Xfg6OdJTkg9YiozhxLVpTmjPqDgahSKV+PZAZOIV2ClRbkUNqov8fHOqOqCstK0
DGnrcde0zpc9/ns5/0Na317yhp7vI7GZaGVCXEB2Eb1r9I1p8vJ1ar1PvLDfOSxNadRHZxFPTbn+
73eQQJAztFtceRGGM8wqmUE3P0JFBCRxXabvSxi/HylF6uvzEkGjrVIEm/C9lqELp8iRFPH5rirn
9QjbUW4vmzu/mDapANHF+rTXe0xzcbFLjpXamoT8T9zmRgH0JxdgNiw3oIAIC7S7kVW9Nzr3tdnD
KrYmH80B14DTx5C36xYtphSRLaZ8XExbmv8UrskhSKRZGYBY5Y5Snn7TtzljlPvIDmFG7/IFqhPO
nA9iF95rIEBoXCnDWMrhf+OHsoAR5DOh3JOCahDIfOry8iZZEjVaY32yRghSFDBnfozuZakmh5tL
wJmpwtMhr0AAnr2oiVzykRSzid3zkJ/8kvrcO0AK38RLp8z5pm2AwGfRlE0k8IQ8NO68qiQXycK3
NSR+wlxvj4nERsG7A+SnOJIL+KURvLDRUNlZVMFn15VWNL4LbzfC/+AqWVuaLZUdRqIzMhz4fW3t
1BWBYTreveLFsH3UeyUWXdb3SEItA1GCO9CgWa2nF26WPQKs8WACKwv0k5mmkqwmokyMtGzHtP/0
WXVbrwD+UVgO0TXDTvxJ3hAE+SAdz7/3CbZCLkV53zcEqUr+cT0ByV06HeQDZSTbY+CpAizfPTnT
iS2ZAcEwsPe6X1oZpu7gscYGe2XlnYc/mNSbCpKn2hF8qN2DMa+Yd8YhXS4L1RQHx4YbXm7eYRii
c8UMiQsKPwTfqf6PcPFKV13m8s+qRkiresdJmNBPga9A1BSiPeAZ7O//vu/uo1TYWOUU6MCpzTmi
PQaeUK6oSAKWsU8xVCebpgjrctYsJuzVamK6cJr8I6hF146k0HODSEagLRWjFqPvRlWyTQXJQWcm
awyhhR6hK+tESF6Z1mcdpFOiFj7QlwY68uJt72Mjn6+CN2vJaYNPt9z1uTy0/5232jZWhyvVcwX/
btjVl8GdG1QzhI6hihkt0KbBSCkx3NkOAXGaYbu9V4BAUBota6mHjGzP4ThciUhk7JPwaYhfvgYE
1zKFKwQpSGHcBgaNX9XhJaKwmrEOOrMaBMLXJuNyCxiDK9tfvpgpaS2kR4KsNfALJo5d5bSMP6ey
corZSOHVATcdQH+yNy8QUEWKG8X+l+9Wgfi6IoJCucBQVfmAli9BqzSF3S7TuQidYr5uLuSCgmo8
aIGX3HQMvy7te9iT2v+nEDbPDPrvfjh8WQasEqwvo+3dsnVtqk8XxAsll4TMwV/V7NfjhEXtnDyP
qWlsIZp8mWkJpPfVXQ1GCoK63llHzl/prYLhm4lAT3dk3O0LGPzDb9re7FXDRw+3g+/xLZb1mnSe
ZYOtllxeWQ54DJnoeXEWfSDzLaxGipR8LXJy+PGS9K4IKbo2HE3Gf/9rzrVRyY1KLjlPuHq88xge
183s+DbqD2HM9i0Ixub62EdkoRjBbmpz7Fn2hBdV0pAIYdkTnwJY4QiNEGUYsSkWrKxlTuj7xOy6
vwo2UbUbrq19bHs/0FXTR7gXN2EjuWEyR2jUQKXJbcM506/nRodG4aAD4QpQZMZ/7N2fM/4Irhts
wSelakdveZdLvzDiqZW/SyXTUSMiEzpf0Ufy8qypzY4PMuNpbQJcrh4bWdYXO5cdMjdVe3Yo2tbg
nfM/ObQIphFpMsBgtm40QCn2bgQqXj9U/UoVr6yzQsuy5+b81jfvZArT+nZA2HftFZUMqcLFbROf
7DW+ZBW+v2dLjes087gyF7CefKrvpX7RGh2Me97MLswqVCyDspm4UB6lf1QzaXPnN6M7lnVzJCTl
b2IiEibNWQM0oIw5nMxiarxm2LRn/G/M2xScYwPugqrRZiZ8cQpLAoYRTTIDc/YxXCcDOK2gBG+f
1npuT/8e+x5EGXzRoY+tGsFYHh/WIjp9Mc5nJ7sXrHUT6TQDl8U8Zpg58hKY4X71Ta8ChyZJT1H/
PgKR8OOd+JPHUa+E2b3c/vPY2xBi7YHJjmplpFcwy2yolPCQgH1X8CfUq1KhGBAM7mC7lZkXwOcc
itvbh5gjgVja0GyJbA76vM/L11FAdoOPVcPEtj+q9cmIrGIbTzQf0TD/wE7FOzGUTb8LortB24bj
VfBrsOiSIwDqNNkmhZN/mMocfiQ/VAo0Cd/lvZTzPMnu9vq5Ykhlh4E4iat9KkDynQ1bhZSQj4Ef
SAykX0xMj3M1dOSECe/H7k+0noTr6DOhxIt7muOU+WLraaYQAE9HIdrnB0Ve/CStWyfuXLxinf4a
ZW55d3aLWn8MYvf3J70jvU1Erbr6M3UjWw/SU7AcGCnLyfwNFTL++fMOoPwHA88o6TpeM/gaxWmK
MFM9FCsiskF1BEZdOi2b14fVF0STDmbGz+b4K5jnI8lzckZuGLN8VOwIq53/romMJ+JFiDohNEkN
TBHlK+FFd6h+nEEGWBCxxgAQxp4HaagnAZ6iPNzhaOdv4GLx9HxdHguwBl+9NU4WgkR4vJ6H7uT9
XqIPhSSFtdlrtn0COMiV2hN6tfXZC+/8NU3ItxMMaQaCZs1plrL7z4qzo4FW4rYQxz55omFsHmzL
98Nc80y8zLOffTGR3uyNm0nsGMCiV2p++q/V0k8FUoPAsAWGWfaN10F5wjW8hFMmr6DnBS9rKn9Y
iPky1oSHeXoEVuA+I1GliYdFENICKlbOSxeM3l3O1ixTdOogrLiaLgdFyd4ICZHT8/GLJUdN6YXU
J/M3vP5HKEDPQqJJCQX5AP8IMOe8a5pF3R6lBS4JqcJg0AfQpNJ+oPA0eW9lKlAO9jZa6ecNx9fh
q5VJAysCxUgs63zaa5wlHw7dyHF5tH+wNBfj8vIN+cAK44zzQvtfiUE024lBCD7v7qShTbXbB2fJ
Af+h1l0+vpv1yahFAxupc7C9dhZrgQqVHVG0Qau6sTUoFjCHuFSehwluaCEKsiBypX+DCMB4Dvki
vwpkS8YaESb8ZbpYsCdyCaMwpokfFOaOELT8MqLjE7CtJ62TF0Hrr+tv99wrHt79/OBHb50kzVbx
fG0kZ1E0NMImiVcHbm7Hh1NbUtlqis0J7j/RChGSYPd0GkYQR2Inks9ElGnxUP4B3462EdYxNURm
ab6Xjp77sUc2YISCv7XsH8vYxD1wZAdoV86jxz/sV80t5TfXApCIburoZi53qpeMdnmGJbYnI3Yj
2yWUgQ6RXLmncpov6hjY2DmqtcgT0jOabIMURWOntQxSdewUBsLG11PCkzlRQH9JsAzxrU7SS1Gg
smQFRheN3Qqv5oNfc/0Jl/q359qz1vASEE0F/sHIvoOK/LzeJLROko5ysFCZJq653tOrgg34rkgx
oXD5t49qHTct4c6cfqOdUPO76OmIXTUndao4flcXJv5mF0ZB7ap4ehEgrx+FDEdubN4ufPx6+L/D
pR8ZEh/+POcFXHJeimGIW0VLKSwFGVrHZ0xFArwiXeHV+W9QJnuX9scC+1Cp0d6tLdmLLFxQUEpR
TNrGM/us7nHBKh6Ca9/V56OaDQlZod3tG4ECAA7JGAxtoFTo9x/XEPeKpzfilb/yZsslt5DUvg1r
I4PC9ZvTQSAsUk1FDv15UkuVtDeR1GRnzW3hJKdNWjznjZNUpH9QQikpcYtnH47d2gPF8ImHtnwf
ugTv81laPaSipWE9sx8hq0xXJYO5Xw3NWeg5Q8JbGCY4XJu0hCTv/kcClr/hD2So1L957VTozmWl
mOoqWU10XFWnEn6LWoOs9qDsQkuThrU88B4y8khBfv+SyTQhNFmZixMizoOhYSfMTsf+fi3BA4T/
nR6T0Igdc0ZRG0wFA3QuPGWuBON2dOiDXyEnDziEcfaqJ0J14D78kMdYcf5lCh8c/AsZfPhe7RXD
q9utnbYkJdYkARnuK75ZFmLYidUO4O++5E2zRKGRfvTc+3lgHUPSbdX+ks6WlFn9beX7SjPVEhp9
nXLoJ74DKa80IswbX6AiJuwZDUcx/dV1kJTOWRMtU+wqna1mRM/20PRy/9Ldq050KZs0s3aacEBh
HD1ALvuXpJHNbi3yeGWV8dOVxhIVKFWOyWdEmLJ+DyQo89ty2s+/0n/60bV2tn3ed59LNhmfzvdr
VCTZAeLAHiUtVLXxO/s/z7FPAFBRVYACFR0jxZZ57UY6QejTlgUZT+WHib6EJ6pohudvro+3AYlf
qTPhETkomsh51XvNrpz9pmVFmbA5fDUehOI1ocHNc8gOCqewZGwdDEgZbEuRUz/eT1b2i5vJDIPj
DEqczb/yVcrbhg6vUfqWf1uYA0Rar/DzBO277PRdDdbDG2jmU/ll8d3lOSGvdVuEltTvNRBTV3xO
DIt3zspNdz3yayOsKfuBhsKw28vgvssVjIiYnwc8bRZCd0eV92QPk9+n2XOPZM6vgzG7vF5/cZ4R
cuIzlnz2IjGKF60JdB0wNEEVom8tEOKpEzLq2kVbz/Po1Ivckl3ENXfjZpOQxzLHodI6A4Dr16bF
8Gxg4qkNy4EKEMDfWFSFsvOxILuU1l80yuXgrJqkj0fNk7eNns1A2EPoU5byqB5lUEprByujTUHs
cQaxgXRDuVxSRraB8JaOK4bKR5iqyvrQu3W3w0H9am0FmeIrGy6X89AlqjVGB00l7d9jLjPIT41L
YuwWXnyPnmbGd/OVKrCknqJFPBuXAvdNoAw01FxYF1j+u6nTTwbZHMUY5IY3lYI8Fp4eGRv5Nq3T
jM5FyRQDSFDOt9COL4taz77ryFcUEioAoOiwFfCkGpYzD+7oyuw7a8QWm9fvmZclXNoBu2MdHXo0
OpLo6NY7ooT6+GxG/6zYvOzK3cU14Mdm6MCiVCxRu0BqSkDLNJAqbEQcLKtQnkhzcC+rNSn7D8uL
tD7TtVUATyylxm8GhmiQXp9mily07cZAlv+3n7UwF2HB4jO1GUNfV298pbcOyTc+fI9U9iJ8VGFh
azdTJiP2Nx5vxYQQL/haflJsL6EvRw8XDH8+gTGg0m5sZ7ZtgRxlIDz8gkuCbsxh+4vJdxsvwDRZ
zdoXsfNoV5wvSOpGp5bJjcNiEwgrLW9U/sI3/vTRXe3bDAjmYE5ZLnBBjKpZyigv432omZKKmuSg
3IRW4SqyIjb2CR6CTpT19vlAA6BCsRy9kAjI5h1pBSfhKKIMODM0fb0kBZbDHyZbkr+4P2alTjkm
dLUrlo1tBhoDC6ysLO0RDziZYyDKBhxJplnEEVZmdtvJOBTOLmH4u3YGiglnuumuKhBJLxGV7G/x
+D2BG++9tOJdWy+RGEoqblCAQhjbkeFZNW2VF5Wvp14WlOS+3tza0qkio2eP7HaLvm0swwuHynxy
eirJ2MZDryNBcinX9jKibO8t5ZowXHGago0G23V1NiaL9pokYZkkcBePJ0v5Hp4wZNU9xc5HRM5p
A3EmgjfYmbkgK/8rlGyzo6fRHt3e7fF4GG2z4wnor3jcw26LKYNri7fWJCgnWYWMIp24teGsvlyv
6MPqvaEI3ndYnMVwVg9v5Q/ebhsD1TT/S+gALWxxjMMHVRuWqCjDx5SyT/rA2kycJjP0/3ldvdD+
EbaJL1tnlMTGFXJQ/7g85BUIEFWb2g79JNG1BtFU5+ii2YIv/AAYKpVAc56oFDfd8RXGNcsD5Cva
05AjVQ/7KoKhbMoYlPHnhlPp52KyZyygIPhJuxTGfDjy83O18JHJ9T1W/b57jV44oh6c4QWSUNZq
YndfPhwz4RUMscGlJlfJYPgL9j2N5h5LPs79U1qRQ52NzZljJtOgReB4n6rZYBXYKAKSR0GCpl0B
EeGCVuXl9VB2UI25Nh28UUIk0mUhAwQDBdO5VQhG8DRgD/zK1oZPHsxuR5Zw8lWsAPP5NT5q1ZU3
OTmVofHAd2/jQjCx4YpGWd7qsYxDY5JtkYdj96uLlu1Al0QeZqCuGC/a1pg5hos1E55YWaV+lb1A
rpLf+RJMsm+ckUvC+7YK3bPnaUBLdNQoicn0QUcYaCCFc359HU/vHfZHrhFMpKUxU3jMhWErNbx5
hvbUqrATbOqGQzUIPerm8gapVzhA4WTHloVV8mCQNyP7HIhIaGOeyVNRBuAZHbTN42MTANDVMnBV
ryla0DKBQBkHlI7GWBWB7kgv8BeEH4dddFwVDXac7BYB9/rkyJzu4gL1bFnq3nH7mOVMVJ4obv38
N6BjAxeFKAX87FHXnaIkLtBwrJTgLeIEwz4HxwMELVnJ6yzmmLWJOcfl3BotwJIszjxWvHmcHvaR
T9CD2oolQtuS1y23JadetBL4QmNcp5hNhAZzYaW1w6ME971Rqd9XfowWuXGjKmQJjXuZ8mbm9rnt
qlC583DOvI9mh+n75W2Hbw9c6Ad4kIKlxmmlMbud1KXrmd9V9rI8FAOnWP6k2XVG7sb8aC7s1Dk6
Rq9vC09xm75IPvLOGTo6g7IEZcOSfDuhzNUuCEe84HCrwWc29xFG2FWyhK181yUKsPSep9PAE1Vz
fRogbzhiyfd69nyg0NfQH7orCk0XnGRpMqFLodncyAwBKwgckbzY5vAoieADPc1Lv2Q1S0wPdum3
6xl4Kq8az/1WwpdonqD7GtR2DTs83oKGxtUd7xcNqN8NtvMQSjm//E6lnDzbxTJNFBmq1o5O38O5
Ahd9DQSYdgyJxou0yJ4JGA8Gyl6WBCLEzNJRXv1f68YIs8bCJQAIq1JE/6fkl9zD95fnza7CPq9O
3ZeLQx7uCIRCexcJXtioZf13fzvjxF3mw2U0GWbY0fV2//UJWuNETcSUTBwelGXO1IrbTcabIMf9
DZVZG5u3A2bDNzAHE8HJp6j0sQ0VO5AxPyAEINdo3QRFfLpAadtefgZ8hGKhYsLVueyQDRUmVMUF
EKpht1SStIjEdw2eToqrd95HZ7xEqKUcMXC6Yg0hDeLKFgRd9FZSwQnqovcNLCULwNS9pAfIuKti
xaSLiYoePqBqoV+6E3FjRTZ+cfHuIOLkrdQROsZm73rDm2U2t2o+ku07mRlRW32dG6lwuMCqoTBr
bG4rz/yvYJA9q+7ogQ3Bdxobmhc+BTnTfktUUbOemNIbsrXx04w7K5ENgOK7MJX02xEiPHKGfPrN
YB9B5jTY023X9ivGyYW7eMju031N1lVRR+/K1JKHZUPSoY/6uIISFLUJdfK9j66nT3rfA6pBP7wx
5xLU6pYyf14X6cUskJxGD41VLQDwPw95J86zcMru7w6ikStAnerILXz6L0wCDNQbDwGet/nZM4Pi
fgv2tydqB9U1phtWJIKquhX3OC/n35Houd+35gpuUQIDfmPBNZOJAlS0z8G7MmRjievayzMhWiHX
JtQ47gh1bz3HGLsxx4cboNXyG5Ukts9NGMT3VwVQCvE/ozpaIhcfNZXEzqXuDYW6s+EMErN6hNfw
0GtASXv14S8dKgz8QnWbTZM2rvLt1T28QeMTvZDazbK6dGMnWv2nDiiCw/ERrPe4pjJ4ZOvHEJCF
+sSp5NuQsWhHb4UvNs1AyA1Ykdrf8R4rXOovmcV9aXgDO4dtxd+kjtE/3+CDhy6QNb6l/3yCI41U
K/QcQbfLRK3WD5iWwXJfn/yjtuqi4IpYiTjRhCVY1MxyQj/DSyBBFw0sLV6IfVyq+/et0/sociEt
7qpTyDC/lfQGM/F1+m38OkzwyH4udMCrzfd5DBnI0eBzK7EDw7u7zm7wwzHF+ZBecLjHZY74etGt
5+zbBvcSBRf9UV7jU/JwweGsPrfWD4XSSm+seqs9ZHaNHBJYkblyXhlfkEMTHXvZ7G6CzTZmbwuv
6luVf37Vdsz0gNadRzghow9S8g6/y5fOPXQGSJ/9mZUiVXLVPhNPPuLviv0vazrY6oEkEP7SdsUU
wqFgU6p1THInaM03H5e6fzlHQIWDBm25h4ItKOkkD6RjRmRGnqn/kzC1EkoDlEFGY45aSlcMvkFN
fOeg3HTjbGKY1KEHa0VaDKJbXrb5/JLojcpOCdtMIJOLeFUUEm+dSTUV1knKM2zDDAON+Ju6LqpX
GsXlkl3reJB4JEYfGHP33OCGHhf9ilhf0zi4foIOGYySj+z35gkRu+4eHn3PZ8tEBIAl/NWs0mPi
c7VSxMWsAkqPTO1tqfQgzrLdg93665ppfO5/3t6CnEr6DMaxLBcHvqMnux7mi/sixOx7TKdGsOzt
1b2V8jc+AKjuBTvIrtJ9e61fY42XSHFDKw1mJ2x5EvJZQ1tw6bFbfmuLM065Rh8NgaHeJCd33e0K
Gn8+uXIZT1ZvIAYTStaCMrmzl4WK1YVC/slGzvySYG8US4V1H73gxttlPPqsVH+kEWMFOa3vk+Ta
DtX0C2crT0ruMhR7lbVl8ebsZlycl2ff3+yNcQj/ZQJlj1nYwCi6O9yPvxJQWZN1GzTV6ICdXsui
sOABKGTDFd+DZnwjqVPu94EIPQCFMzc9B38MonZ9iuC7sBgRuXGABbqGhMNNKTP8hzB7LOSc9/M9
C3hJCRMxCXtZ+YbY/FcGYYXUm7HIYIgF4IK6zku1ncWFC//10XKpKySbXxwKSjwkPaypcObQuOpC
FTpXdfzsB5OxC/L9yVMIk6p9jge6S22IIZJE4h6UX77n1IHo8UVm34y+VXhzd4OVs1PBbbZk7PHT
4D5KBBuQ++muLzCp8wvy/mJL6yyYW55VzB6ir6xwGxh6nzwP7fnWAcicNL/2OTFtBD13T9xI04D+
w6TOxpo9IC75ONvl2oHkTtwFFtfVX7wRce1VpRe134AFm+9tURrsDXnDdyMi6fOMVNz6bO+ey2rW
XtQVdk5jy5RaOsV6jedh6MRfixLi3nihklnPqNdYxlcDB6rhSeaxEdNaqkpcv4LKssvgyyk+M+vn
P+LUIzDwWJcLDWwEn6rCXSTlq3N+pjTuVbeGrWjdNWb3uhSYir7ey0trJvXpSG7Gvlel8sPiex7/
l7CAectekf79KeOUD4LciwZ1aDBu4W4uDnzeLUlBgX3WkX35rfbkLy/4EAmdD/Glfuoq6mQeV0tv
TddNf5ts4pQnDRPaerKzM/YKQ1lrAiAowl9QGua44mnK/RPvUHObKGaW22fpR1nUtbOWLldJzjqs
ySiiA6xKjG7RhgxKOt395yWz576H26BcNgkwnCVnxC6JrwVJGitTBpiXCCtP7jpODcDLXV/Hiw8n
NWcBVP5GggLao/BjqV+8+ZYn0k93bxLxPEN0WFIrZiYesoMiRVDvgfPwmuANbRLS61F3CS7cBfdu
l+Hwx97ERj6tujytwSiIqk/JBH54BrhH14M+juqK5BBEIcgsMVTES2RwRr0WOh9BFKCdxd/zHWqr
hYB83JpkdeGuDOvzH+9X4+R0WGLIaD9JjhcR9F9yyPKq9tpttYkEZoPbGJgFX3uaYZ07tRWrTbhN
iGpcKZgrDfyWMF32tgMltAc/FGa/SC0GPo2EoDdEJtm9tt+w94mbQJHEvXcTo6sn8YmH18Lv2/RL
KNKL9JoLGR0JbVV+lSTxJsc37bSvhz6Xbm7iqhMibu2/a9H9CxcFQaC8RvRNnexyh8CxxzpGNolX
XUMP7PENgC7JYoFgPGyKlrKw5UOvgrd78FTs3c27y/iowlvK+mto1x5pkoKz5RwxWs4z81+yJufX
mmzhF0PCse+F08vZ37v+Pjg+qqCEBTkSreUmFM/I8Q5lUnw4N/hMkhJj3yFgTPRzBZA1VGEcx5TS
Y4YNhU/mVZv0GE0mm8ZqUIi7QveiW62QWLu67q/NwyzXnteoPLAQhh06f0aK5G53t9hDAQc1AWxf
MUHVGdIjf4cJBVHXcNgh+PWvLOmwtJJLzeGgBqqgZFZDAF+2iUYySUvN74k25a0VxncEgSj+M3N1
i654RXwHzf+roF4W31MYpaSl8yYfFSKMPD1mb2LcXK9UJiSPsPahECmq2eAfVe+SxDVN2SvMoes1
LsbGonNts5VvuheIpBFkY7ci0tQLg0poIO6WsAWdSlG75sD2LrlOMGMtewX6d3eEl4SjSlV3RVvI
kVqtEn6ua9FCPNW2/oveLfUKoF1mWDGsrPu+px3UXpCtTy9rvPZQiQbywluTHrvhbP0Y7wKM9FsW
OjSXULGKMsv4zFnOfpfwUEXzAPDBcIaqmjqqE+M+JepuxxQ2HDtTIGlK1LaOyTm/3USbDRAQi6fz
cjP3XfCN8FmqMJ53ik7JDGqYDHqrgkahmUxmPnGxd0Yjm+PDDMQKGDnvfVVlBtJZcDat3C1T9iy3
ji3Q6HwE9bs62blJCMUsgK8dxErTIk0wazyuGL/gvIOyPraUr2Nv+kcFnBDqJBEsoKntZOYBrY6e
c30ntWArVnWAZWT9K0pSLILPKeIHK7Vmq23le+ewD9XCK6HePch2qpDyWQDvi6Dg19MSQr1p/W+q
b8fPioh1xSJHYO6y6NOirz5hpHk4UqPAacvJ+t3xBwCVA+CBlPBCFhVpNSIKbTxCqG/KxI5a+QKU
lLH2ATr6914/VRu/IOjdKfHo9VC8y8OodBao8skb/3ZKOML93DGvE6Y8oWG6kC638sH7wTbBE4Eg
cReZXNA/Pg9AoiuDtBMo2G+Ye2M9yGKFrlsJn3C0tNo80eSNIqfGH+wtxdVQmnDAdY3rvDBl418c
wUGBK1iyLdikEZ3fWF73GDmJxKJPEFmTI1OnKhSMq86/1MXcRH4J0qmPxjLEiPnR8nC6B3ti8/bm
H7KEyf8rbgJdPOCHrNOtTkcNa+FoIiHQqYDlID88cR5qyHhINR6Ku3yq/7ZH+nxilg1kgB+6+Y2A
1PAJDw6Ri9AdjaG9drFoMKHwH0acA38U2/672ewj0zFYb+q0g0n/ysZkcSXQ+k1sV0TMhHG48R33
MQrzk5TIRf4N2NNPNZvryW/asb6IXZBGDCubLHLPxz5y9rAnMH/ywohDMCsCbr42rouzsC7W22mR
eMwcP6jQDLXl8FhIk7ZAAeS7YLuus30eJYR8dnN/9BcUTcsVOh0fDCNMCC4bDTK1Kp7+1mFsLAFZ
8Qg4g8OQoUbxhzcDlY8Ej7neaBgATqMs2ZCRgKCAoPqh1QiXTS8sLloyKoDIKAi/w22LafEZguyN
rbgOWnW8coLKPj5xsnr/0xIMvqZDPkNTg6/R6wSFprDwrYaYKU2zFtXGx1/JCKthwBsuso9RdZrP
rT4xlnOLBTOItZ/Yyb23xgVQ9iTzfhsEr4gpW3+njuNzYAHGOcldO2ys7IREjByKZ4dQD94+Q1HC
Rs7HJjSXy1dsf51J1n68Yx/qD1p6RbnFSyfGHQrZU8abL1j+Utyz9vINuRv0UAJWc9Evi36FL+84
M5eSk2J2T17s2Cb2LFtswarjswTmhT5IdBvpSwojzCK5kIbhUymkglofEXrLBgdz7ABxpH9ewE0J
NdpPy7s1jkkhVPniRm0amg6K7Yoz7MaRJGBYOBpSAs6rx9IEyJ8mgvYGk0+481YmKzV+dePJD9Dy
9WL15tK369bN9uElqjCwPawfk81ViB5VsD0ZJsTjBJuCj9aqrF7AZK1ouMV9OICBz2WYAUklPjS9
YeIz48dv5kQNjcKi3uadAx+0muIyxIzLjN+26CS50V5uemXNxa5VALg2wc898wp6pCmATi9YUjUq
m25rgI/FQPFGjNBgSRKXh+rxmrLBEXa6au2GzjLCTDWiVtF8z29qAdXnirckI9Z0Ifk4aXKhp3Be
Th5d4GSXzGojOPlogO2d7nUj7qMO/q5M6yqNuYsW6RWgjEiWfcQNArHQymeTrkBUrTFhYhOvGNt/
+23R17X5sNUIpbvGs/R6eiPpoTdKBzXhvTS3hsohV9YKWt/tyhJxDLujUZp3tSo0JD1vNYKmJuTa
g+S7G5GP47xyLz3BeNxH6AQ7Rjk00X3ShuGJc6dTSR/Gs+lQjia0f2HS0JHVuW6vSfPOtmPYnSY8
5aJpUfo9tkk7gIuryx13E1Vc0Jd6jFwluLgPF0baN8eLAmkJwyMel3b5gHrAtvWjlK2ZyDNWNQyb
3eccs3UkxMHNHIbPsVXSV/lKNsNruqz9sRSlnGG738ynXFRT8YmPcHKKQNMAaw8xqbtzlpuHXR0y
2b3xcRc9z1vdpEk+NkItdLLxiew+E5r4kQIHcOv7YP8srjsT1qynE1wk7LFiatpIWZIwlS6JjllV
36MahgPGMPW03gJR53+ZrxLyK0w5wx5vBgjV05A5KwEw83uZdkWo00kr0pdyBCGzC1OnCdJlf2fn
+9A+Yxi4Ap3OX9Jx5kDTQYcqPRcSPkTPVeEvrOYARMlcSgHSXWmTG3j9cYDiWp89+/MyTje7UMZO
N2JbBcEke3KRVvi33AI1gLiCk5yw1ETgi4szJplAdbzVAHSs2Rey5wRrXhTVpEws++DTe/xx5AfL
AnoY8eUPMMtY0UmXkRO3ygBpe52fYuFttyyWSkM+7Zas+NXDMUdWcF9c1onjooxb1ENwip5p82iB
I3KFPKCIuLtdeCyT6G5eql4nhB+5nMHuy/gLhjGOTRuHBv4cGfNwMDYPD4IMa1OIH7OoqZim0mAI
xXiBDP1E1qzNzg/bqgmMaI/uMmp144gpHU56S4c8+pSMUkWhQrL9Wp5TcoaliGOJqiShuq6OoUcd
Gvqv4uf/sAkjYzLFF1K0ajQp4KaN+CTSseg96/s5XaWYlRX/PzN3RCGbbfZ21cAM66/oVO3D517I
lHfqp+RrVoqeoooD/yGnP7AY4Dhs0nkLpxCcZW79VFSX0o+zQ8JS8hxqAbvLWimzvKaAg4eY8Psp
HuyES/Qk7hb6Z9wa+31RTMuwZ/RjwaStzYa6a9dBgZjsnHX9hQ4w4vwcCgP9uGF7ilX8AriqSF2N
TymRpWb8KreA2i0s6gAw3ff5hQxE95sMCu57rg8jxn94doDRTBuifeM5Sj4s4D0xZ/0LVzhSA+Ph
aJdhyVEzXGugfzv0iTx9ZbB7l7o/1qmuBIsw+D5Qat0N+0t1ipYxY1XEJrwFUh5WrG4v4KorSN1j
CO847GpTSUmWdu4D07abTJH9ewwudmk5ben/3zJ9gmVA/Axa+0uXO8xeWJmy4zCRKMcrg3h1ClNQ
P00CfPchyVAu7TqajDT0SgvrpLQRoVPuQ21+2HPGrOWVPnGgWGwuceKWROxmVDdXdEa3K/s20HW0
9SxJAVDTvRLUboqv1PIhJQRawHgZYNJPjWCx9yu9gDma8P3FICxsAXIgTTQIutbkrrOOwMbjSGlU
ZoQ8nDGvnvBONn3o651wkJCzUZiyiaTgLJxlu69xDM8IdNJu7MimPe+E9SSqrow+/oDUp14Yo5Z6
0KMOeNPGENW6CHAamvoMww2b/sXlU6j+xsSGAwaw9PA/035ivUjzR6P+K2LTZON5jXCTd9P5RsIu
zcXNX0az7Dsiimn9mOL89H48ALAE0npv0iYBydiLXW5EqxBpWvzzPLe5tVqWMv0uQSXBoTzVEzJG
ATDMNekAkbC6hLi7SHygarQvgS4ejTi3Mp6TqutSpxxWY5IO6bG+a6G3E4in3iIjJZg/gMH27klh
z8Ne3XJ3VyWS1hPmzBs3+qpQ2rdgS/nCDwS9BSo3CqX31qd3qj1iqvMEp5puW9Zs8I2s52dTDuiE
dES6RTOiPBwxvcUq6WG5cgvdwXeFzUrOepkRWbvZvTg31vduTEMODvYU6cOtIX9ESF3Ew6g9q58X
h3gKnaxxDiCNHlRoru9XpR3yl+CTk7iEUDGRFujoydiMFlVwXHyb35Mm1WC6vtDuDHY5qNgX/Nii
orIsGKfBBJoykwGrlk65xjDiw9LWUqOimO9DUIrll4Bz/b7rcas1SQufg6hnf8HK9uc2naAu0FKy
pN2SVRWl8BfPP9jeCutcr4tdRjn3+ldagSK2tuJct5tbDtPXWU65wbML/PKTUI75te46mtsweG7Q
6qJ7GKcgcFm+7GwABPqlkDzkc90DOtv4Q72RG0IDu5WpGRjDAGK+RUKULUGCnGUDPXuh2wAEem7z
ODXwAST4ReX9lg7mqq2hbk/EPPmx3c8auMQ9hxMEI67pcs33JeOoLsqOZa9i2JOYCwNZgida2D+D
I3NNqn66Tkkrfa99PL+RsfhmK1da2Z4kQrrbfTLKVtYQbD/cwX5gQ+vH4P8WH0gUEIzdZFxZ0mJx
B/COIhfNANNJ/N7qBT3iXp0mg//dwoFNUTJkDX7R68fG812Oy1H9O3tOCIvBi8TE6An2i92mYjB+
2acOuThqlZ4fON//AahVlMYzOBCs9oc/DU2jFgTVqACd0fLkWf2bA8GvfT5wdonLd0U6Zz2hBgzO
cv8+Swxg8BQanGyQN6valX9f9yu5T77zQLS3gFj/NEbQ+ZcK3OulVqRg5b8OmyCVmi6gwZ5N2S+P
ycp8mSOd0TOfME2wFM0vh1x5RhsRX21vaagzoE4TL1VK9+FwphT4/EguwG4LhUIaAOLnrmnBwLvT
v2H3I+6VowYQ3JchOi5m0h26WMRb8t4ncPhdECzRtMPo+ZJlp5ZdVxvC/g64Pvah8ENUxJv03DJy
+PAFoor05j5QWP9Ngs7MbeNmgveTCzhhMNuc6Sgbc7ZAF3HJMik+3xM7UVyKeuTn8eDgBGwd3QPq
DoUMPvYPqFb5hGGpkgudrhb3CexvtjkqXv48ro9t3X3vXKYoDBIi4SvnuTrCxCtQAt19zPmUY/4r
xhTvZ46EaKArDlbtdpFunIqMv8VkQWJVmRwRMylBZHoG5Wv1XKJOmdtIIPIfUaVjMBrxlSlqQbDz
X4ocCy2R1GIWhH7Rn5EYQ+FArrQn5tTojN0KIiuq/zZ5jE9cnm1+jt6sq89YCN4ySl+2El8AdeDh
VF9yYMv/0sgnuNGDlCBH1oaaykckHc3famOF9Gwr+Yi3YX1LFg6AWz45AOvTxPULPEpYghr3A+7S
BwItI2tz0P7+Q2V6GdjndZoFi8DAe3GAuZNzyKO6Ydq+oAVRhxo78rHgxxcBXj8wV+HeeJ7+YHbn
qrxkhGiVi8wIJ14cRW/bTLJ/wncRD+suolHL5wRKFQx1LpDuX8BGPzygnTJWRRQl3wcXmqr6OztB
mebuXuXSd+6YpaP2su1EE5j2JR7vzBB3jVv9n/CA37J77nA7yQTL8eU6JlMaL3p1OE5wdtVpNfBg
M2PmHkXgiPOh6DtWrR/U0DDeRO2NVtP26Z8N3R7OGnFcr2U2rvidhjMxLYONTpA/fVjCTUFJsVYK
EyVvmIDBQvfCTM9BcvafuPh/8EaJEg15D2M2ARpf9+OXOdeZuik50XSUgnLAswDKwIlrmEhlD6FT
Rx/JXmj9+qEXFOCfdWC0cVMbSyU7ytIKpb4KbVdEnRh97HA03KVRukmF7Zd9OyV7HNYV2vmWbMqY
UWKBafjYEsYy0bTwcf4C1yoNfuU4p/n/UwDEYiGRRYmXnTGvpzxCgGXZs/GuGAjctJrJtvdzzcXp
qNsjlpXw/xGRX5UfpXSb0C46yUg3EghAyE0mdbPj3n8wFZQ2Fj+JqolqVSw2Gg/EIzl3tggGnfLX
hO5kACkYaRnBibEq+Y5rlN3LcTAkcHsrRqimgqdeq28xvexqBdz5YNO80ZasOPndcBS0KgAQNyTf
PrcqvuFNfYxZgDIDqL0wxyzdP/D8FuuY8DmM6s/Pm/qjlvs7CEV3EGJsVsLpuRa8S82+zkUxVAJV
zh/TUAC7MeC+S0LhB24jCJiJfgUMLiFegQBC28jbe8YmK6EwcwXkDik432MuDj3mijE+AT4Vfnxq
fUydqTSx6da9a0cP3+G7A951vFxjzM/sHF3JJr8yD4lmXj+LPsAaHUqE5Zruz9lrJCiJJu3EZQzO
WAMKkkX4cVwA0KIJKvED8g66t5dqss/NGzopaI5geCNhZd3fxMw9+qn2f7HIB/VaZKcpfJt35mFd
7AQ+pYhLEo8/mS/ctfPdRP6pjAcpM6m9vMzyIH/qo1zmUCf1TMXJsB2LV6D1K/kT7NAOLOUUJ7/G
P/7LWskuiN3cN/6tzZEy1GewbOm/1hu8NCPDxXkfxLCEfgzEVZxUa4SKSanHDg7IJqucsnsjELuK
dwZPTMi67xEErir7FvGZMGl0gysMHjTraf8tuutEi6Eg0CtgPd7b+7tLoDqM2QG8BsNz+g4a2I0Y
Ux5yRjO9JlT0PVnrv5Amu58anyOopoZYuX2InKivDKJr+kQxJQqcmbyEwVOi9vtoCv9DU988Qw8y
GjDyNUXWKw0+ygWSK2P6j99r16cgWk/Y9SJjWDFucaZZbWHDfA0eem9VEcZYuyDF2D2cn1HeMR9w
bTnEx+m4oPMkWhNym0Jf+VeRva+Z/6wOmDtn4yyrvDZySEIxQJtZQAPtVALOhubCYakJARxH6c+g
z2uxEO1SUJwjW/gsvh7o3gwGlz3Fihm0A9a+msYx/FrKdTWbZsRVfzFFk+O2WGHBKOcPgEt8FTyU
0uoamsV3JKWpQdeDirXpQZ+0gKS4Erg5eQivYluH08xhj1NlsNNT7b3MzkKykh6ux7HAp32ZPaXX
ytPp6lApDBWZzIHEg9kLfLvFLMGD2grgCj3c3a+rXqTWCYH75B1B5Z2ibfGFVtTzt6AbKlUX4gVs
e7XPK2BQupUjqb//P5aREvop+rEusKNsvNiX034ous6YbOtPy+gOyfsMRUhaUXYLy5ee8kCNUWFG
c0+Hez2xKW+GpEP99JImUq0ftBlhseeBWvauIR0yOKq1OUbxTWMohmjLG9VshjQIXbm6d4l8ebYz
xP6iSlho6OYhLEoonn0LM2ox+7IS0EBq4FhooWuiRQq5G1RQP9mClgbRFvA4eBCXCNax1aGlSDoz
M2w9Kn2fq1GYsgpEN42TZeRljqDl9FO5N07POS+pWnWaRW9Wm1k9gcz7ZYPI4Vqwd2YVs36nqnPA
0PDpWNmW8NeFOCiFkBiFnbh44FEby8PsoMZblKBQWTaktsyCKAfkCA7bQc18hPmUVeHi/M7/X+JM
bMOODZF38wQjTVZNBT3Ttkd4KsoX0WlvkjToCopjivGYnC/lHFVUbN8He/8m7daJG6qzY6nFn68l
wohCKuHJGNFqOiWUJ72vqtQkei8ZaY77eSnXsaJgw4vBOUp0TQyCsi8DaqE2C4UpdyOWfwYWXrby
bu1g8nsZ7Mt4iCIgCsDeTHHMF+S+XwO2+ksKpRsHuPdvu+3Kch1i3MWSAshYkvYpn4XuYVZw/+Km
IAFm2Hi7iB5i8ckVEkh12/woeNw1ZMhpHqSLfGPz9icaMcOQCTTCF4K1GSRqOaYwbM1W8nC5Afm9
L1mzCX9MRAoK3JmhLiaNOFgJhmkAuKYSmokhFqwAc1WjrcnDFsfGTCAX8RCX2Q6jytbHIdgLSGXc
pVkKN+AGQSdMSeN1EH3of/ldaJ4n+NVrrY6AREF8sTL5izJPrOZXjiAMpUrVJ6hMZLg2x9wSahFU
ZkbbR89HdVszhuuboPr1CGCFMrXtxfpFvA3YfOGcgiVSpUxF2JOghVrSDdI8w5YHvpHuFMbEgi15
4wK4aNp/QayUujJhUldchex06MO/xBu7vDtP/VjTKSPzKCGS/xPO6kz9fv9YrdH52zULDynzoIqh
05l2xz6+LqDVTftSwkceomNTaNICn36tf+Imk/S8y8et3PlQxbVTHNIoe4ZpDyBKuTtJRLXTKAAc
SGiuTzMDYGCGcBmvwWoNP4knkzUC9pr3Zsfi0PWxCpUcKEySDEgDg46nt8eX8T4KdCXGXquYCSsm
RIic1kQ6RzYU8zWiLDu9RZ+kGHQx+mbz5lxt2Elj3TACnYUc1XaPK6+whWqzAb2TrvqxScvX2WJp
cTlGLzofWw9h7R+SUqJJWJYKrZ/O5bhaFK0zPQqEDqLQJzdh1y7oFybpeXz9WPSm102GXCCYVVOZ
Aa3Bi2071RF0gi7xBF+8uEuKVqeGnacl+D+/GoCy8h7xLi3l8oPgCSzklMBNN0pQlHs2zccLNscY
DqFiRpWF6O1yu7CcOs5n+/EYFRfc3kd27DVCgN5/3pyGQ56Vc/nHZcXPzbo0wjVTzEjHsBPb9nhS
Z1sAfcGQSfX4qaUDkhSekXfKMCwZ986m+ms/DyD6k0uPITMIrndz9B8ZljLt4FDpBOhWyKBNjtl3
sPyy3eMxOs2A8384GxAQnDL5L7TtCutXEJ9Y4X7ax0K0M3Y/hZUFIEjEXXRWbZVLrGEUKiis9ph7
j/i1qBv9iWv3Hbb12b1T3ywHc1SMOy+N7ZjEPSRUnEWc4lH42904XfsVokvWltmJ6monM1eiyD2M
88z5/61zErMlOIVYpA6Opkb/xHqhzEErx+ZiTIgKyA/ow0YWHrzgaDer2w1Fl8BJOXQ3Orfjq03i
C/VHhWOrFPJsGoMr320bbu6s5cxcq90loWReoBrKJFdn83ggfph6InsdB3Mv0NBdF8KLdmbqZw9+
5VOVWT5os6l6mnb+Y1Huz1oziBsZ8mZR2Xnph2lOOmH2/sxtMjop05KdOPBN+uS/hy5S1IKb05qo
dbZATwZUzwxW677wMbKvQrGVzP0aplkfRc2PY8OfsZv/2XNAlL2NNAXpyQs5gO7t4V07kJu4V5LR
dxe/cLIfcjn+QQmH8mLu2FSvYfL940FWFGqqlF2OSaAeDXHKV7EhM3EjaUortcDaRmuwZGmg0fID
p9hcbtNlMX5Lf/DACkx1CFI/J9vHl6mB2OFJUr0OVzjGIQyXMlg1YE0kHET9CT7O3z6I8e+h1US7
vFl4OUm05NSNqFheOkm8DRzXfUzOd1MYortalHf/34welJuwx9xYNVWY7TqJnT0lS8NgJAc7Qm7A
3GrcH3YjN5iZo8l/MhG35L92Ai2XXSARezLIWxmYqQIhPZUdBxI9IALv1GKDwcVoKVwxkU66ACQR
m5LEELRyIv3nnSdojgmr5vmGzelPTkeueXB7uG7A5K8G7VwtCaXsRuKKknWxauzsAstOX6M2ERk3
0JWLMKuSLCYWYKVQjfdiKpaEPzCWx5x4rKKZWRMmpaz3yy9jj/93TkVaRG+kBq8PvhL52fQ9KrzJ
Pd96dlrX4ARkm25YkXt0fOcX+FEadys3EHv3RDRcL1iY8NStnz9JGCLl1ge069V5974GDu6OzD2n
71G4xJXQ/rIWBic7owZ+KPGtXyLWJkEC4+JrECVaZ/YwH2GemERZhx131u02A4VU4c5hTePn3UpK
XCHglH/0H0nQBsTC8HLIBam/wRKlJeWucAIL7nn8U7WJKWP8ohM0cB1SFUztwxBEoJ5CcnmdsECZ
cyp9uvirQujf1u8ztG3O1wv/O1o0zswF321XhSpLZ5Snx939Z93YAbyWQ8ERV6+A2Es7VUTkUB+A
AzO8pdNrI3TE1cvvw/P2To8UvziLOy6kQc5rSt0qjteT0QeR5+zkvmOt4lDC/R1122oA87Zslt7p
BEPlqg9GYpHRKNVP5rUcWHOCBrWrTbhmOA/o+2ka9csqtfxBQrMUqXKInVJkQ9+YZyEOofTyAuuV
R6xJimXQMtVz0qK+nTFkjlX8P00W2tQAzjU7i4STyUwBe8cPGqB3lmHOYW6ZeOglZtiMHxcWEBSD
m1+ZA+nTTx9W/EP606IoyK2XDwhEa/93dKNpHKt79Ps8S05rRFUX+8iyu3dNx+e2DYPzYhtZJkeS
tpUPU3NKWKEo1XaN8Irycoin0D/gqCx1eIA8jcIEtSZ0naB98kvkU3+l03kZPgHnj6sRiNAeFqgm
R8ZCAFek7yD5H4h4S4oyI9rEncmq2f0AXWh+ngVWXbxUuHckvVGwr2jn+zBjLists4SU/QmXY5V6
oz9gRLM81r6rzzF6QnUky6AgrPQHCrNwO75YqCxd4cudxCUpoFY86dFHdxVmsW/qnUJAaPCMV0FZ
GQ7k5bBpVh+6Am0SrYDAmEAqutwLEZFcKwfQYXWG6aVY6UeMg+wqj65WY1OAs1uEcd8m/RSmQr2x
Tdwql3AbbhjzBTvs69QwHlW48RUmsqrP1q+B/dYeti2ia041+/D5XplkZdGUOa9I7XrTwOl3PmvK
4N9TkK0h4bC0yQMTRRUVWjUUNjlBzHywMFVS5sDb7C6ZBoOCsIq9Ks0qaYOfRzWIzlcBkwnHMpEu
MPgtuYy/6P7H28c5z2EsN0A1dSPxW9dBi8sacI3V8ZquYDC1KocpDU3HaR7sCi9YrHXPWjiYGa4l
QEB4Zsc+mEd98mxC/B2mNmMVTM2TxnCJoFZutXIwtkieURYyS2mbxR5ADLNHwARKHXwBHKeFmNyP
o72ZsOGkKVIpBPDCCXhmv2kc4j43Yh4mIVzF7Tz/KwuOrSzS6fOWD4CLSes5506jOkufODSPEeda
ggZpo1B80b0i1Gq2ZC90y/HmqED/6cc7d/m/z163MJt1gdNInke3zonURADRxMkkjLJyE6fYPqjw
NQUbRmNdNQm77bQBkG04pannhWudW+f1gXMg5VS2iKITLXRpZG2kYBBenSMvKxvEeyyMbWIxWP82
uOse4RbwuH4Oth3jAune2I1i0dIgmJtpTCYamwvjXTo0sjPVz/wu+NNaR/V+8RgsojYuuGRBe/Ux
C6S85dwthgRHdVgFVgZ18JQk1tC7YdgdozvYLppeexqcG7ggcb5/ZuH/o7qN2r4H1hwUcbmKEBxF
gnmv82NLLX9tevf/PNqxZ6/eeBipSBaWDmIH94zh71A2PwGfQIxLGscBQu2ECaL+PBXlUsPhv2YH
MCY/o1fUYfbogstbRb/kbpBpn+aqB6KhJLhIFBTeg/B9Nc171WLy4Wg+JG02XyBSnGxMW9cx5isI
RiD4uerbaD+xlOACgO9T3RI09+iLdzZazyC7tfl70+dwx8lfpu6MrfpZi/107uvpkvT8cHS9Ui4t
ja4sRvU0+FHYNR+0qcmONekpMSAjvbJr1Kqzuv1wSlwr6VcAER9jwN5x5Ju732BhZ/8pbis9DXpx
x96g+KC0NlRJk/l/BKg6zfnhqsy7KDszTvgkjUCtIdkX6pMt3E1j5DGdTxSWrEpbOQQtcSl32T9N
j/83RxmWzKa/L/TYPxr1or6anZ1G1f8AuawXrRL+MQh3zNdzGk8nyTjvvUW4JXiNYqcX1bbkTAil
5uHz06a29gA84Pf+PRmOj+7KBJsZFcdsmEfFQdul2klLF7sZkkW1sp5KQR4+775UYzpAxnaPAKWV
JejP5mBi8cT91uDobVlxv77TUTPG3Q+aWF5Snzc7yyjvpvpkmxxFDVU6JV6qac2Agn9kWxdBGOLw
rrqrfFejxEA3oVvbjiIywu782idTTo3IeO0aUXkjasTPwny8WYpS4+J5mZVgapydB9oqetpHD0/6
evJ+HvAaoFC+Grtj9gzQqJJ6716PtT0uC0oD8+gz/yJtnMAn3EwVWKtb9Q99GSrAtyRSuAIzJpTS
guUoBDFvplBVYk1uBXEXmb9pwv0UZXfaKOrcEkGog/t8kx259xWBHSqiw8nS/GyzOP4vOBYzPuqu
QBFDlvUoLCSzRE+oB3GVcAzUTRLQfT0fFhlMguHusZYBTjhcqvjOU9qH/C+4oBOvrFEM4NSllg+O
9dx9C6Mvnlpxu+RYnFJoIpV+L0x4tHqFODLi/COa3qvCdkgnmMbczXtsUjDvdnnlDeN/qHVWE4sm
T1cVu/FJYdH0JCfPpvNHgpYDNROJEjDwk2JOCUvCXc7VC8mP4m4agZjjbMeRTuiTRoILDv44Dtm6
75+NwTZJVX8AbHU53G1lhlVRQvHEeHfReAPOJ6xh2JS82GzIxQaxEweGAwxXXvSCqg6wzmE4bkVB
Sa2mHMwuJhOQJ7626zttT3RBUoj/X204mhJJeuNIcuPU2jAe+U+pbuxGvChVa2HfTdcWgrMyn5pN
RasAYMdt7TgS/2he9Je2FNZy9oV5KVNg+iMYABfTVsudLbw5/44gah+OV2jQ0VhNLjeG9PPhmziT
5Ywdb0r/jIypLiEuM20aXhAZ6c+2stmEPI6Tk+AWYefdXJlhQ1CknZFnU0oOBVjAIaOR3gf2CSxQ
61vmIyKg0BuB75/jMPMojltAx/EnmqKTNN7K0bOM7k5EHdlZJ5wo8Q0JW3QX2f0ZssQMck3QNs5+
+5nF54SEuIxIfKzKzLrTrnUIsI/RucnrTDDIafiKQa4ltppScxl94A7G9d0qeBBaxzWO2xQ0SkKp
5izo/6k2ZBn/ivk8qtWA1HFq6elPwzvMEvTEs1t9/2Gkby6GntRC+VgFdVoihjJ5w5CTLAcHHTiM
qMVYagidEBqCfHDVwXHJHRUg6fAUxkV+jOqQRBiE5D/8bl+ADmko/n+Jkne2dK3SP/7FRckpC7Ty
/Hu6dQ3+JmAB7iTfBKt2TKcVuvTG1ZMiYq7pfm5BBYwpYPXr+Tuz95A6wyfeKDo8Mz3F8yxQmIHa
+f6pMe0m0ZXxIzxPFlv38gW2EZM1Bl7AdEeKv0C40sHERD3XeALW+4Q5Wx5tJzsuC2gH5AGmna9C
lDomgQTQJ/bioFQZXHGRwL9y6tworwo/dw2MTBPv6acXKtdWtremiJhKvEjsUrxu0Mtj+y0rZpFq
ZGGP4xmSRbFSpJSrtAmwgH3m263Vcl6lsSm8Rp70JWIYSk8hOwCoXAVTopH6T3rj5Q3Ua8H8BX2r
E87dzc0JE+rdpfU+N1w7GuL32OfCUdGIszIIrI0uQWq5TPFNpj95snj9vD5ZQ2oanY5EWJbnG7rO
CaQKhlbz+IXkmhhMqNCM85PIkLEHec7uzL+GBJfZJfI1k8j/HWtZEACeJRDLE0bHzg61GoZy3UW9
ajK1XaoynXyMvZbwjTOWWnogXGJ+P4W3KERONusqqka6RpnUzn6D5JISoc+ZwhwVgibrXjqZRYHB
eKkLMDBzzXkxRB6y5mLH6KFGaSSJPPgvZKfWRmfbgEvWD0tEjf/Ngn4ZOu3S27gmSBQEcfqdWofn
BVvav8JXiezXcmlyzWHeb1KtBw1EfOU5peDlan2suxYzRA1IjwJm9denJKMe92d37pnIxBgctPdQ
fMp8eyYDwG3Xrq8JQtCSPvZfjgMTqF0L7MmjY/3rOsycwsS3bqYP3mBOhus1u4a+IoLD1miJB7ax
HZ95leaYR1kopHs0ufaD6O8s0KCa0qnAKSFfxZoLdK+pUnyfKMqlAqSlX+KbJTz7TTV8S0KGXLLA
h6vxJJiSi1zvWLIHWz54gwczba2SdoXTjxlXdpjfC2rY7HxL622/tCYhFkWeGyWwKdnEuUdFUeXI
uxWqCQrPzxJtPRYshRDyR/UoSufqck5ahw1ODDho77/ba3LtiP8FhhJLZiY+aw2s8Zft9kdGU5Yw
RnJEKBJLmzuZ9WNwtrulaC08Hprr89NkaEpXaCatx6FmNVYIJ9NjCDjZXgMQ02+H8b1gy0Fg/vRC
7jKW6X2dW32r9I6HBjwGeitYv/cKXSCxcfirdpX0jwFNZgGP/HOvQdChplKCDs9Z7B++wQhKPaS3
1/JAbm10tRqjNSSHcOUInAkQXHORUw0uYBn8QReu3YOe9ZHLuJcsaTfD7HjaangQgFU2sldyuRXD
/QYzWCD1QaDEsRknjc1Zg/kVp8iR2ZakkjW25P107HgnzCvpgoQBwoccRiB2v9GtCZymwNT4SwU/
rnwM7ebPfnH1xNry61mzZ43MdMc38j0KmG12l853+GIy3U3/zVy4V9EK+H2oaXSQd/6ayHluBvVF
9ylF6iSKQND5+1cpNgsawn/ienXT7fK5l0ObkzvDvL/iAcM9eN5RcozIPowBos5/j03QVUXiUpco
M9Fyn87f4U+V4AK2qHep9qunvQSAQBnvyFTs9pdQLIX7X5so6Of/TTQLWxaA2QKC1JBRLne+kQxN
lutLBQlVW7tVj9uE6c4c01ofcBm57YcWek9CeYxQ8A9vwWBUWP3bFI5hbYCg3nD+iMsGymFE7NHv
/bGxhHfdHNi0YEyhWEGraceObERcwNnNoMYJR0HRRn46fctZuTOl7KJ1DwUTDv8u522tdfK/2Oxp
0Xn117CfXqADYHPlaC+r62Shpr8rEGCMqpmrr0VMFrvkDb1FzMqTU0CgvYHF16144N7knJRaXa3T
kJ3NNFVlZAcEqb8XF+3g8XhUOxGTEv1I059zHDOQGZvHzP3WQi0O+QyvjVRSG69jfUoOUoqGEiyr
U+9rF3Zz7w+GhWoyN+jYODMmtrhzy5fHtYLeb+tpHUhe0bzDc45ADAH5cPMxXo1nPI9LOSHAJyox
pMO5u9h4cqHy4Kt1IRpqrJ+aJ7QW5rIeEZfQe7GCosbkHV48N079INlhLnueuQob+xDdG/JB/REv
m0WJHOAKbc5b6Jaw7w3Ie0OFfj1PQF8i3RyE/tkU/ZYF82r5xDuZJIAwSIi6eCbyfsev0fqhX10G
U2KU9FHJtsF6v6wLnFT6zW+BsFaA/KxRsB38trkJ0h0OEqRE39r/pBQCUTNCxN5/pE1oQAcqM0Cc
BJGN1s8yg6m5SPK7DHw6/lSkNKliCM/EiF12fvcxJzi23krwAMjiFAuDr3Z/5gkYTZ3UD0o7C3Rj
NFhA65Pti17xPflmGPhHT3UgWvW2UAhZMLplVW7rNktQ8vAMjdbxVWnSApV5eZRDSxZ3nqSb+jJv
VIV3YJyeZ75Esq5MG85bhugSd/5Ldhy18ziTI6yeGYQIirkg+dMKZ1YkVKt59xQiDf98A2WQh7p0
X1PUkr42Fff/D63IteHha5LUTb+sRVXg/6vK6rbQVsK/OFxNiTxdra0J6LGwVYMFanJisIxCsT2f
qIjWXznd8JLqKA7ZWKgs+n3kN+i/uD4qw/nIg2V+Sw0RyRbwHMwFr0JuFp0wNnC8Mb6qjKKrHPRg
UiqlDXdJFi55V5/V7WJBm7lYTlbzQSdJ19Zl9xnGQu/eHR0xITWh34AE7xPSPP/7wx5HUG/C4zsz
FzfmWsfBheE0OFtaTg4bTiSXQ53EdDBdAvEc+AyLglYExS2xXAPs4zodHmX/6pY912gfxPpPkxXn
w0SkbUbZJEmcl1RY3jrY5nm5DkhM6ytKDnGAccl+FZAgPEqTKFxgxK28WCbGYzb4Ai9myNpDJwNh
F39LNqu0XAcl0K27xsAW76i2uzml9v5Rqbmsth9FEx5Ftm6gmOdye52AIWOUkHyJYYF4iTQwv9ow
iTUmdE26YswZOtNyiMRmm+M4QvKLGrpnCxjEW47bmrZMdgZRBkMVXY8ghfuZzLLaGeSRmStO0htS
q1V8ukD6c/O7oBcPCJ0KQtmHOjQMsfsJGSDDnLg17vaDQ+JeD+zJEqLCOuxlLwirpv7yprM2SivH
zzUlnLfqOfiMnpnh0SvZY59vaNtXoimLBzEwgUm1LzfmufDaC9S6JH7739WUuuGFp96oDV5okP9B
PudTyowuB4CphrKxC93U7Ii4wi/p4njP4cGH2bgKn4TZcXQOMgFGkIFoP7dOzC9gEAxBOlH8XGkf
2+GYagMj8M4T1b6td3urH/ffuccuB7iw8+34CsHofYOqzq+7SByuI0RjnWBsRC0zeilPYhyeswup
1PVmIZJmy2fhU1aAjz0CAIiFK102bJMcLLAJtUlogUp66IbE6DTxZYFZ3LuyOZyQtZ1xbvpv3aEJ
mp0e8Bpnlz7hm8JyyZtskf4CJPgQw3mLT/1Zr8BwiGN992gRzg8CFXihzyyhekBChIO0UUR82obx
FuZPNh2qnwnsJFIASEXm756LKr6tRj9swFUanamdEXkZ3KLJpdDSSwb/uBlIm8Q0Z2uuP6gtfwwC
pfIYVQa/Y+6CEBDm2jMe84vFTSvr65JX9gWbalVlWMo3cjZv+iFiUfLiVd907uofWzmUipNaoIUO
K48EJf5BMgxO4AEsltxnIv/lf6B8AArNSJnLtokRy1LkJWBBtzOazUaX/UkF3Qckj1urpYNeTDlx
axEywy5HV8c3NIObSSXHrE6jW/KqbUaSAoONkJimjM+dPTHq203kjtUubZotbfdTw7ByYjCMcaJL
8XqAZxMlAQcxJEyxF3Nc2F1HeV3/NlG11z4YsbmGYG6kUM2KaBD8295vtnjylDl4C4DOCCAOCGra
sLUg2qwgIVgVOfyLd7GDV537H+gfoI6wnmV5y+jfDSw9Hul11IPEE5ziksTHjU4BDl1dk89v6iqa
nnrkVUEcjcu7pedLxvPkus9gubkZgwkWCkI/zehkj42ETvQL4Zvc0WenDdgMZuHWtpFw0O5LwL9Y
SlSXO4h2c53XepJzp+x5JFLBR0kteP7dHb+f5NlsOJteoSmisj416VklyBLH8NCJNyg3Z3u53uPw
iqRRNEeoahp35Ly4ScYGeeZlcpo2tgOy8ZHNB1PrQusDalIPjKY0gvxM757SmbAt6sJKDi7tk5+V
tMZab4X3II5Xi05TsNzG7xzypfdaRnQ1tbLmBO2bPsGKpHEz1EqG5kVLIFk/T4lxY55iQT9IR0q4
F52u7YuG+IyLlNo2eWf0DoAeXTCBsYRbM90P4ZLWLIxzB3Bv+SAujMXTcHZzzypE6LhZ6LzQ1PlZ
lqraUdnNhyJeJIdEcbCV3oIfSNj5CujT9SP+Px3PgZ0qCLKioI8M1v240wK9CA066KS/Akt0M/M9
gDYM5r6wL6B+Xz6HkhDFo3ezW/fGlo0/XIqJi3ULzC+GGuqL77nwqsror/f7IYDGqeIs7YYFFI3K
xoWuZF5g7Fa7hgAlDIsWQxNT3zd7MyW3iKoyNI1xmkVGxbcCDHFuFfICzK3al6i57KRK3knC7xXW
LQfT2GILYzgT0Aocf9Abn6qX8Wc7dh5Aq0uLDbrzsxa9xk3fz6yHBLzxfixYuPOMyN6+4e1wDxR0
Zay4HqwJOC3D2ARNntRH4rZ2lRh8GyQNX5cO2RFJjdq6ZCRYPO5DJ+x8Secml0ReMaIfZ0WAA5FZ
Nt+EXf2GR6g1CE+j/tgDDfToUb7VU855m01UTj9eP3IwqbhubucurTQ5T3Jp2tQbn+CB7yDHoRyj
fqERlJlvNrriTcg6uuAD9ySYlkrWlXF05B9+hIlWa0jBVuC7IzVjCe+XvyYzpIE7N1mNy/wNpKSm
MAKyk2h8lGY7yv2gkB5/MLlG1Cyligz6AlUdv0Xd6wNxIOLuZIbjSslpWRoGkGBUCRBuLRWQp+yG
+9Qb13Ax1WiJvQh+yDZsktHC/JQ1iS0GyhwXWRhitrbWYDH9dS9uq8Ja0zeah78wXX/LK+/a9tzR
8UPS+lQ0eoRJPYk73m48d3GOedAnHGs5CO4oGp+k5EPzfY3ear349TCGMCkbtL/61L5SCwhHn/oH
jCciRmiQBmlQsUqaeDC96CLpq5C4fhi7vKEzXVXVe+2HXc9K0MhbCF0RwnzWeOaqTB2zvk8i1WH3
jYacPz3dQMQzqnMOwjk74dB0CogjwimlnDcmE7uIL20NxlUACJBmvd/T/z+FfvZ+VLSY3RRFcOQk
7+EkNi0SLQK3CoDeO33HLg/TIdo8rW33XCFtGIbcWQ/3sM1+NEKtaYL/QR45ai0L169ryvVDRioM
wsFDYEb8xHQ+chD3tr6etahoSJ+mtWfRU+ZGh61aAZFhP7j2mX6PYah9PuhbFoqNvWTAsWVCzsXW
WvxtZAhbBOG1QSZdOkghlXTD4zX2Yb9DSgy/sQiKRmgtcT3VcjRo2mxUlqEKf8nh9Hmd5n/dBpJH
YQF/hU+0o+9+ZXPbM4YsVOWUaZuLYcSoQWaNBvprNHlp9uRP3gcASw4HBWlG4OuGk9VkZI4HNBeM
5BP0YMMhnM+eEFbTZ9cUbKwKJMFgd7eiREqWn5vJ9Ehg2hNQ2uw1wu9tpd1bsTLUknxBxl63nkDM
4D+VH285m8DHu10Jh9tBTOnnfMztzNlV03WAbVrET1SREuSVNLMK5GldI4YnDBI1mZGcrAP2GvTE
tQxtIr9nRJKnTnUuTUQWDRoxWhf5N+t/K3zQv9iyJUGATMZS+/+jdE+XWjlXdxyXzHvmwzgL7MkS
ISFeiHSkhaA4pfN3IOANvzGJedNppEC/sKv2wzlkd5PZ5fkjmK+5aOyVgv6vVZh365DfBYMK8BxP
hKGMkKxAKjWcCkjri0E598qnTxPtNisrkEjqIOorr0vrZQg4+SpkM1ucJQBWYsCEozE0ed1sxiiE
poHlMSUF84TAMtI4p0PUJVfVorjZntwS6TDhLPQj7U/DwtSHVnB4vneru7VReehZ2bBFWfOzK8FM
I1xZebFiI6waNRHxJ3K1gcdQi4iKr0+yYOu73/U6nJDbkGSRKzw0ONEQKh9pMvfBv5oAbH+tgcTJ
fYNA4e/vnYpWUDwIphQZtnxBIS4TZ0yuFuTqbYZG9Xp7zc/cZv9GMnlC6G3MmiWF9w5MS931L7hi
B18dVaeOS46eX5FfAgUzkXXN/KJ/1TEIbZzgiS6lh4a4xYpnJoX+gnStZ9yTLeierY+u1SaNLQWL
hzp7aOBxZR2+usSBrRbJ3BhpvLaoPrD2d+eQUj2rysPw2lZO9lC5q7heHRcdJuXs10NLq3k2pOwk
QkR2whwBBVW6406pXTl/lEPxwlc9IE0SctF1VKefvrGhFX3eKGzXpS9MMNss1QWP1D0kCac5+Tnn
1k4ffqiTjsd2pWaspw50v/Zha32PON6/Z9s8+IPmZY7ZKJthrf1Tc0ewWrM5rrJ3elwT7862BncJ
ZTDVSjrT0hU0q8Rc/ut2QOMlSkw07rWdJCzdTss0qzybE/RhYFSARBMAPCx3n+jS2pdogqI78+g/
gUQLCI+Gi39n3S65EQrw9GBilO0iXGNwoCrL9n9t2LWBDNR275qt6A/WnerMlZGuAHl6aHTu6RoF
eLoHOwZFbqt0pH6LspdSBMRNP4oQZHnhAQ277Ql+O8pCbmiTP/24eUCZniUS8wcp7t+kXA5eKPur
F5ljkxROf/4c5jb0EJw7b86dRWeon92TSLq7hxZACc9syVc68wKBeuHQWke/6tYElsoGk2hgxT6N
DqxWuySnWexG5fNksXyc+XjzNo90CR/urijXHCJnpdLaphf15RdvJlVdx0h209HeqiI9mOti5nR2
lJ2/uLMuXPDTdQREC6sSDJ2HzfW3No72fAGA1Y+BaeboxFkq5/XxV+n7hga6jbXBttRvKnS2Q02p
9yY+ZXbspc69rC1UGIUh4fKlwkYELaFMstkmApguf3mUse+S6HjOyZDExjozSncKn8GPsmQhU9v8
lCtvIvd2ylIjGnUw8e5kehbMxka5QRFb7JPqCB0SzaIsnc/w6Pqvq/ptD10ggmJRAiMxeFCZtgaN
Hr4blqFEic1wLvaAFr+/VJ+MsudjImpkFm592l0EKSJHvk4oJgH+14u97ptFaR96J1piyclgWFTR
ICU74fgDR+9loQutMUdfcxu5PyiWgUp5AgOgWaT2yLZqNmywTSl1tTijRktxDQeP8SVlPXQ/6mD+
d9FebSzlXl9drPkyyvPaRX5iWKXvSnGgEiRUNwoFVtWMy5pFAGJuQ6IBmBJ3a0HQi/1wemW4CYnW
P5v/R3rG1hEWbnZ0OCxw5Q9gucT1YezYW68oJgVUOoWoF7uyhflyexhoNkwRZjqDrEGokGZYSTPI
DTOuBf45fdLtN3MR/Vdx3UhGPqnPAbS8OHiLVCngjqfI20yVrQHT4J0Ct8U7XS+lE9GSG7grd9xk
0XXia9UQpVIbblYUrz8lK00mXik2JGVNClcWHu+dH9yWTn7pRoN34fI6D45QAbhGSSd+lFPyWYSp
IwtDWTn8kvf0a0PWXSLEJpDY4PaD6CMfpw4Cn8S5wlhBN1HMbKlzcLrY4e2QTPI4DVG+G4STCBKy
oYiV6Nbp9Uk48vBQ0b3KBVZlj4xTXTv/rBewsULrK+7Fpif6LGWXqIZml8Qolrp5bOlAtN+k62Az
3EISBR+RArTT5vU+f/C9hbdB3FChqL253iXasQtZUQ8CxcI53SSAY7fnV3ficY1PVWt7jknRFJNA
71UN+stC8IeckMCNXEDqepFAmzx6J0FVns3OlKtq/L2WHhNNrqb+VyEWiEcrcfyU0fIIWv/HPM5U
kpsJ+1iLAHzBFzNrScVOHVECnuvUNTBe2dmv/c2g4hTLeFtXB5qcwlsJJT+86vKUtdFZEpL1BPll
EISOGsesFSBS8VWdeqU6W79l+1+gZ2Z56PF1Ui0VmICqHfwD1FJvAEgiKiFxV4U7wxhz3kfiz135
jC4R0MqnhCVbDEZbbQ22U6+StR+Otgxsvga7SJEzpnXLd4riRG0FB6zv34u9IaYIh6pInS9w8Hbn
sZOS4wn1JKDCCO04PgrADz9uOSvyQ+RNBx/JDy3b+KE977iUrLNWPIroOaDUE5G7AieNGFYSLwG0
Uy93wPLGMgIuc0vPQvKBngOzAoOezt6cPnZSMUuITivAmY1wsFR+Yrupd1QMuKmojdZZL+IoHdjq
WKCaqTZ1g8bR7vtZsjaF1UehItojRgV8XdJhyfFPtKHgfmWQakmAIRaiE+sGmqpQePwkvEfVz2uU
evO1r1va8QIWNzLfG4gcR+DIfnQyNY7sp+csIu8xFai3QhpY540zm+8wwW5grU79NjZMX9iY5+TO
RN3gBbX4h1rKEatP0TeShu5bAuqEke2krWpX1EyA+Dc9KtRGqqXhp65Zjq+vkmbOgacZ2wX1lTEe
G21r0AJsTkGk9n9yzPOJLEY/l5gcERETi+IsN8GeA/iEzTYoifDBf8wUQ0jSlGkdrHWT2dMCtnwN
8BTdpPZyjKBIm0C0lAUoqg8oiOASKqbrj/YbLOcBEjTlcWDWwYKxfELuXiXW8AVLslCzjtOZxSiF
aGbTrEijN9VCUkl/WkYoM2tGwHoEZjykX9x2qETS9te/9qWB8phDFXLFMy0/fnPmZZjgwjB7dZen
o6ToE1+GL4p2ilGQEYVCNHFvGApJXwbGht4w4dRMb5vNEaxX5UBqhWANkY9KdtNT8TdRd0tqSeDv
FoTTb+jpHAHF4gQP0G1EBmntntCvW0H1sevKCkofNBTAJaFPhs0Qoc7FgGvLOxUc1EldvIPRBHCH
yy0VKvCqNn4LP2tEJkw0gO6J0yWzOYNUUIVG5iRVlNQVdHHPkdy0l0NbIrDv8F9mblckjzrPfP3K
fgXGXnJ8ystxXoz9SOXxNY2rZ5zfQaqe3F5G4pHDMujZCIHnTpbm0piWriytVIIw+ORpgGcNG+96
VVhN7o1pSEt8OiR24UW9t320w6s/NXu1tT78kINI53CuuUxuVP/ubQbZd717uR1v08KY1qhSBRYL
kKNA6KbSIvDhZ4sJ5h55rYOkWqHrnZAP8GI3Gz0ZWPW9P9dIeegse1DKSEzgnC3WTxAv8iVqHVhp
lgtCveq6YdkYmvmRcFQb1RfkXV9en3UAvkZvBUQFYwPdF7tZrjDgPqrxii6Kj9J+4Xn50xeZQ9ox
lkI/rfiO8/4DCzxfeQBjsxNo9qdEAS36B8yG8QFxUe7QRTHqaUjqqi4Wyi6X4ZwZDQEuIEQPSNoG
e56/q/OhrA3d7nHHrQhywgEfB4OI5s8bRM0dUMjWSVVyinNTo8TfamX30aEpemCwaPj2CI8VMP2e
OPpb29HdrBCPLaKKyxCUhaYO6Qlh4IWtJajNLWaazBerqwL8IsryCy1aeDZdq/7Rwfh6kmMhTr7o
+44o8f2E1PlsI+7EAe5NzAyqNmOu8OKh4o6buVFAmzentrFIkRI3/UInkzuSxeEQ1raUgVAVRZs7
iZR/SSWj6T4m1EM45KFk4Xo2V3+LWk2TF97GAyciFjJh+b6MFWMeJgqdwehUSIgmz7nwuxImV+J6
2TCDgk/FYMapZ0E33s7YdBkXUYYByDxyd4CjroJOA7mDPQdcY/S0qmJZQiM1LRF5CMflEPEUJ3hU
3EZ82k1N1ZeXTEddE+w2ezE1yOFg00dcz89H+b8h95WyUJy6Iu1PyEnydrSPlKBRibZZNxU4VI7f
L2q+Gci174nPXcRXnMlU4uxl7jZ0L7Dnbvw42H/+amxBzNKW7q1bkSA9qZKZC7Xf9W3yBN5vwGeB
E5rCLj5+sD7XlNSVjer4xw3h/swr01q5B4uprb8RrbdZW2X7RZgS/vRGwy2RnY3y2fbotmTfyPeA
gfEg2R8Sxwc/9EvCrlJUqoOe9XwBv25TxtLf+GtRtaUkM934x9E59OJKPBrbSZ6fgB3Qa1BdnNVB
HASofUGMYoi1b13YFL8EUIlxgdnBuQKQdB5VIBXrdwEYnqWOGJmkwhlPtECmzruXt1kCiNRDLBP7
+ixu4PKYcEqGJGwG5A8LICeV/Fg9E5nENkgF9mhqPLfdabht+ZNZFZC/KhNLcBZgpl39obpMLA+8
gcQ+uGOnlxXajZALrZbOwn7zjlGDAt16kYkbqYH4n03+aNNfFcUooQ8E/FUeeH/+vJbM5vC66RfE
6arak5NhlLluReK8GDZJlDWtsDcG4zUDNQzF7bBxDfUjr1UDLOUJR+2T1KpYu8zTfASN7RqxnhfN
mg75xr3kYSxI7m842EDvfH6NwrJYzx74EWBh8hrJgptrmEQiwbGij2Y1M0jXIVAJQgkRyRf/vmox
Md7hVM1MKG+tWTcmS5dqZzpB3oDb2QFs4OSvcJjmxx434LES9lldf9sSWL12zCiVj1KYz2SvC6Vl
dypT1CcM/MQ2hycpeC7QZmdTc8ADV/tzo4JL9D2YQ726MvBEIdQcF/omMstOnqq9554TFPPztK6i
kaRUUMbWJVYRswpMu2JkV2dSnpS72I3y28CqPEf2Aivt7Sr95BcmUn2KDm3KWE65PuxKBDyzQvKT
WFYXI4TYuWvI3RgJdNv59LgOcwjFLh2A0vluIqgq2qKCeiIs5u4fSUaZNY+UP1Iz4tNq7RCD4VaD
nmr0PBkVGwzRxW52HxI4wZJVnOqrjZr1OBG6IvXHsdtGmjIFTcNOMXlmaGJKFWnsCvQVVdzAqoWo
6GQZ5bwgIj21PRsp8m+QC7Cz3+boLZjLbd7PMB9Vz6gFUTk3wj101yC3l35nkJC7waZICee3dugJ
VD5uAaTXfwPEB8Uky85CT7xlrOUfFbaY18GXewkDz2FWdCX9gOSThclmmL/g3t2hHx2YAx9HJ9aO
0p9YYxCYOhH90Zux1IHeiy+9kZJhQ+qnaQozEfvHWRKcP2AariA4uc+3o11kePW38ikVJ2XRn7pe
vq9EWV46GfgTUrT0irvX5lIuNqIvT8DKVx5O0Nb9Rw6ofdxJK7kuxtR3ZsMP1YZ8kynmctYU2LCL
TxuTz1zDi/FuzqCKt5lq8FDbUyjW38BTxYUjg4Wh686YqOd60Kdy7FXRyoFFmARDvKkU4xPQL5+Z
YYPQGixSHnT1ea/8iBoKw8LcS1O8NhIG22z/ENCZKnOX0ynDSy0YJzLdXNGc+dKzH4XQ++UzzCVg
Ylqdgp0R1UftJzlH5sks1grwJZfONKd2EYKq+ftjQupWGORl160hRBry0UkI/z9Zn9cq7zzuRypA
CrtS92nu4maOmoCbv2RtunWRhUtdV262PdBirULChadD1X4c2ftPXHw3YpRShBFWMGWGJVFHM3QG
suqE9O5+Tb+aBVnBt7SGLrfiSaFbTOkilhCS2bS7NAElkZ6sXJg0P4j/ACq+Yt91MrOszGMCGDvh
mJqCOJP/Y0MdJjlYKTkynYCZbNwtrUimYUKfPQ4WJwdCsdaaqfI7UwXmo98LoeY9O++RbjXR5amu
EcIVzBUOgTyZmyC8Ym0fv1EZKF+WCaTmIp1NopVf+w0HpKY0KjlY35YfohY1iykgGSPhLGx/mvHm
stHamvl8YD7UmOIDRR4gqoGXpFnLCoJK0w3zNplpGFBSs09FpUnnmMNrxK1lALqQIKt2tH5xjX+i
o6m0Ch0Www65aXIEcVeg2+ZslJ+n1AZzFjuZlCcGhw7EH8WQ7/MMBxjL5bxtohb8fgPu4CzSsXqh
xwog/HJ+p+tGxq6B7QOqp7Yn8k1Y9GDenTwMu7mwTn/JI9WieJgGOdjfLX+80VpUnLuKjo6CgQ7v
GrASbnty5DXNnbI25B3FpTISGxDz4y0yW0AuqfwiJ2cqT3q/mgi6I1v+eMYlIGXX1yKhrSaPlF9r
tAtWgCQNtJfTWsGbFIwvBLn1ZkayPhrEeDyCBlb7um+dI69iR2hkkAvhmp9Z7522MddiQOgE0sOL
rN/pFt/CKavzkczv3x4cfbW84JfTNhCQTkufDGzgONZoZ9uyHcJWDbuThtesqsnMTUQLO+QRrjI2
4ZQtGS9aEP6vjoO1c+12qnqcNQQP0BON/U38EnM1oxcK7d6w720FqLCTO38KdHVajbROvypl+02k
hJFjEiSVOY6cOAHLH1NFG0A6C82e3kTVKwHBYxMO8Ae1+AQTT6Ub9r5vJAEEgUw+RcqlXKnMLRs7
5K74OUc6Xq8yaT+vuAgb0nIQU/emGyWTGzOpbEabxCsepUG+JkLkqDRqzm7HSg28XalKcwypCPu2
vxYfUvvg6bzGF9qFNNr3KF6QzaaRySPj7wgavjl8loKoB2vbcwPLPwdVEfIj1HpYjypKE69YVhO7
1zVMUvEvduOGBIj1SBshZkwAmgHrg/LcLdUpE/7yU0yE2A5ZZX6koJ7pxcaUlH5yYlfyWxtWlI3b
3FilqKu7P7Os/t2MwNBmcott85kOWwDgU6dE315efk7xARuN3jIjyt12j6+KUN0SEdN6BIRvrSyf
U/SwXdEKGSZoIApzguSejqwW/Hjvjfw8sLrlrpWRvFx9EMDmdhBdcNu408pOpKtTiT5BpSlBNlTg
4zfelOZW8c0wNXUuUu/RjnswnXo4WXsQQ9dcIBoLqiCdxQ4rncqxR1pgWTH9p1FBmlqlN4VzDD9a
v8OozBrhNjm9aAR2qeevYrePEyyFmnO79ry0S0iY+AaLmUO23Qu0D/fpiRQEIKDZu7tFRolqAkmC
h6nSXNzpeCxj1+8DsK33Tf3pAmMaalMzOxsDypiUy/CeN87GHlNymyJierNSXV3IbZI4lK02s4Fq
niMb1wVOiSwUPA6huIQx21wlMP4jVWWEFJOz7CFY38S/chEk6nfQmGByTUO1J27f+KpSyF83CpaF
a/CrtIQ5TtSzzDeLlcEIelFH0oimPPj11enqEZEZEKgXEyegKOC47ShY3b+QCGsFIm7HcJakn13d
A0lh4lc7uPFCOioWcU46737jNNwgxaAJGwhWEyT/mkVE2ZQDGKJP8V6LgXMvNWFnHcX4SFmwVzuu
zCn9v3TDx61hVYMKInJkFL5P5rXfk5jE1WsHygxR8l70i6ayrxt00zb0nnloRjSg2Kn/qMbo/DSk
/q4mbse0zkGzRHyi3QDnb53o21msmOr4AuUOdJ2NOXXB9q+BatQUidVfjg3wH/RNBHFPrVfNdN6p
hcUaN7bjXw6poYyKi60SUU53gWZZqUdVOXoACG1yhGA/PThYlDs4eovgWRnoeKCBGjDqO4CuPmG6
8ATVcCJyi31NHIdY1NYmV02R/2TYY81NptbZ8ICIMC5RV41fky5HI/GgSfr6jw9Ak2CTN37o4zmg
Mgj//0gV/2N06d4BMs0zi2WsBVpv6bjdIFVf5XDML9iTRdq26u5VEUx3FWaCBCtAFmXtvD98ALCa
DdXmmDhfMVRchYbWqOW3LTZuWnFPJ3mhGjKitWGWlzi1X5ENrf8KLSAR2Ovn52wRodogB6Ve/cNH
iF683s5Gjw+tHzvNO9XUStOTBsYXM8rcL5qaSucdK5Q6PE4ZFoMWYGB0jM1z2B/PvEDt8caDYClX
FrQTDXBECtjagTuh845pnLTfRordfSMdyURegHJw9knLaMWI1vAgjJnKHrrdZsnp9l/rC/PwPAig
yH2QdIFK/UPpkJozj27DuEzSPoZl6+rLnfWCgHfbvuXWIxum8YdiVqSI3eWo0l4gh2tH1LfyT+5s
lIPxfjAvsfvJsSlvMUx+9rPwZ/FQHGz7aJWFrsZJiIwxck1O/z5hFtsRGzA0MXHTd849vj71UsDF
jyIqrdlxmtfMSN1ji8/alSZd3V9DB7CvxFFn/MLa9ro99MCeW96Zzaj20rItTGkPY7g8+T7O8ufT
Th4t5Jhb4I/1sHj+Y3ATpun/ti/6rJLnOfw9SGYQUCPMfkhdUbBTiEbBt+xpe01PKb7T925FDOOI
FWL/Pz+cMS4mwZKkXBU6iQYPqR2umKmTAVrgFltn1xdzkKTJmHW4TkSxyGgqzcVO42sVHuvxBqRr
wLXDMVKGc3TQ1CXzklGOpNIKciZhgS4dVBYmxm1yt2tUhBbWGZCsRdkKf8y1p1RIPUqElBhsAVd0
fwg8+nGsGZVvvivS52H+zH2mc41RZBUgnkAVOHPg8ASuGjOZS2BZE0g5xyEb6roRD4Y0bn8QGKgt
p1hi+LCSdQENBSnCIKt+XETSKOojCD5JL6HQJvmi/iRNGIZfmnFWU/JzsLAZPjQkjhmlmMg7UjSp
BhCNjuTpqTPkcspLhKblTIRtRZnWHbOk/DTv6t5tp4AW+8jHsf6f3kYQFX4/UnFEgMKT+856HvM8
AZY4ks9UUikWX93VPlEwUhmqa1Z9rgVly4395gSjhx/qEuhwOdf1TxHesxN3Y8xB9ojy0w9rvF0N
01SGoKT9Hr7SCZP44e55aWEg5xl0qw7pwKejnFomZ2J/mQ7K37bmvefWY0qcabo9yW9RqdQaf9FU
LcjbA9cmkSJoWoPmQKAm1WBvT4elikleafzomDHrEMncsar0oTrlFTl0hunfCi8l7XrjR5+N/qqB
NSFKY8+JWb/plsefRAPktEuy3fFtOSiVu6xswehWZQyHaRxkKV97qacssehU0P0jWkGooCL1QBPl
UFrWGkTRdbX1ttVaxZWmYvUFPRjnVvuGvWHjL4WUAcSM8lWkZ3qvPM9d2mEl81nqSOvsRpdtjd5x
cwivqzwI4rdjennnJp7/27qMvUFOJu8jNwqfT7w+atj2F1+unO7l9BPIqacuuTrZMacdxT29A7Rj
elh6jFjhRkSu71PDVk51AeDS45O83BoWemicfTOeKBmsBQzZoqDXEsGsfZHV4AdDkGLBR/EfS6Pv
ar1SCirHbWQR4lghVUd7/F5R4EEBdDa3+dKQKo9sRhSylIZbrdNEmkjSpYyGFvncW8vyCWVERL4h
2oIPLXmIPLzXtyNcwl4bmGyweiYWZmF6AweO+eYkYHytmB2cKtM8Uv2PQ/teFHFMW6QlHL32IqNQ
LjVhL7aop7OY00ngV2w+Yv+zEgqqksIUi4oHZc4Fj4730QhGa0bb26Ro5VLr54sRwGlc71p5r+kn
KjYXbTF//MBZwdnFm0vlwNlQd2u25lH+xGi+QjkqZZjj7+uL9lOAz9p0cW+Jmfb64GVfzDJgdKfO
QiDjrJPZ2LyNYwlUuF/Gda074NELSK0xJ4ifSXJKlXQb9tGTBoA5OoDkNrPchWzz5t5XOVvNCiS6
B+yDDJ720REoFkqjbTUhErNoUyiB7IjQysFURoV4cAFI3JmEUqGnvgj9eXiqJCQhI/SWZWpJ6aQf
JF9GBSBgQyS8Dai1Mg9dYxwyjUxy9WOqk1bhkYKy8+s68q3U/CAW6d9Z58y9tNiMrvv/9/5oCogW
ruWHrlskksSvMAi4/hz/FCDlmvdTfaoB++a7N73JvAbgyGG5PhvXYT2MQ0eAB4AFkJrNG08jbpFC
rts5zIXpBdf8179n/Rdk09jSfwq0tgNnTnpAq6rSo+d4p7eRCYguYDtn4yxtpIG6Woxu9WrApFQ7
ULo7kHlypBItbz45ii4EyhMy31IonR2vYxUzhf+NtLmrN9j4KUNz3YTABgcV9Uq8Vmr+4X+qH+1A
B70xCpy2rrpCQ06oheQtj7lGyMvdUHPejcdAluOcRXrhOGSFEKpBmqBJXmTNxY3I5cca1KNNN9pq
k1DtSEKHOyeQ6iahkkSLFMqMu4uXIyUjATu7iCVDgHVi2bKaIZLBIm6r9E+GBbDz8OYcOa1M/a0i
JRTV1PY3yvAZ8hKGyZ6GVvdBKPxmncxMZJqvKbiPJ9UP4Z12rkkd7ylgYFYedGamRcWzZfuFJooa
acuvzGObW92gQGdmc9JxnBShgGNdIojYL8SOnko8J2qpYsNSoGaG7mB5MWUnkILf3noMRV3freTM
hUHfcONN1dUiJNDFEw5BvHI1I44MP6WV5ZU0ykj6JawrxTeMX6e4OX9fTNvZMkv3gRVa+FU99AB0
LlU050kgYQ0M91lNviftZe25xQjIJyx81z0mkghVP04+f0dPcYjkKKa2g0TehbCksv8lUtbHmNaQ
dzpzd4OCz5vS6N/SYS+Tz3oQdZGrQI2838MiugilFUO0Kd0dJ0HMiPGcf6sxLsqFryX8Ma7ivTko
kHm1BlrQta8pEBo7SshghAKNwor4EaMrbmT1ggLoeCAd/vqNlC6E+asTobE5HJAnH/3ErBH5JB7G
9ck6jRcpalffPboNaoitDyqvDddtGVILfse6L/w4lwkaPemp9Pt1l+uYa1o7VbPKxE+jsy9f65dN
UmvhRl83p8n6tD1bXSISFmbPSW3VdGsWraFZky6/0VptlEBebwfTsPjxNdfhWpuP3YniV99xhdxY
8cdeQ7W/j5WBUarZO0Ky3V86nc5sLafeLjqIPO/1YMIGNBgmjNlpbe1gEPIH7YMjJ8T7LpoIglrk
YSJoUyYqBDy+K12IbsMKXfY6BId+c50llpoFGRRP/RX4wd82g9AW7ysUZ3z4XaGj2WJiH35FXYgh
Sq6EhE9M70BIHB4t4XPvBwwnkJDNkBnWTheW6/mHo+s5WW0hKXwOvMNtLOibOrGs4dUVoZ57JKN3
vU70GI9sCThhgdP40LEKwCEUxjh/JCPx2HnFHV0EVfpw/IZVgLZb06S0L0uKZ3V0dR6VNoqaIqbw
zOyDBnMKTuLjVHZP4L3XZXTn2R467cmUb1Bo8BWgzsjiEicTn7wJst/28FgtwRJpTltVb4u5Uvr/
3w3Mu2hpN8ZTIYEteqKzkEjJB81h0nTzdkbjpXlj76vP1/45A64TQWU/5Wav/PRFfcsh8aep3Q0m
XzFdYB9WpCQP09hGvucEkIOqyGa2eDxYu7LtrNj+Y7OPKinz0A5MNsmmRFlrScXhbjXmG8NCTrB7
VyDgyJwFzFHK4obfd3g3WmSQ662uy3kDfNC5O2063bEdG+2Nc2AipTW1jzp+SL+8fQoYuEzQXv1R
ejLzJhpgPJyU+naCniacjXx/zVZze7piP4ZQyPR30fSSZfvigyr2eB2Wo6TQaRsR65P6q63IS4dA
+a5YrL57L8heBmPahUvDiWZdjz/HTJwBzh69TflzrF8v+sSsuVxdkjbGt7YaW6qeIQnrfbjCUBAL
UKCIysvJ5OmRu2gFrVWzOHomjKQcoonzmkw1Isxt3vW0xDaAQMuyHSFeskOR+Vypnihofy+R7BNe
Z3AwJac/jQNvoqkfJCGwCWrb3LPqRBsyg7YPsI+fwBBPfl4Y5/PuY0y5kENIk8uXfsyi12oK371o
s6O6hTxGRWkwKy4RcG7Ce7IEHY0Tow+dXPD2pXKGcpCnhrUMdihgDU/nLe/okN4RXND/GfuFJFO3
JuB0lVXqNlPo/aeIsedbBUvoBpf5U9aL5S1c6reCzKu/+dEUFbjpR7+b78Wbl79s27/fDgFI9FWl
nzS1MVz8KX8I87pcCFShxZUbhvLS+RT8MlZarEo1H/T90Tsx8dwKG2cnqWss9gu4akpkq2Bxf1pb
YRNadtdL/cF1EdEf16iPNqcLQrQfKiu8nR4UJ7CKehLkHzUOE39bckXmV0GWO0dg0xFhAaCJMn8z
MOXIsAEtKerhkBxxx//UznLapWFZYY1PQPPzNkNJAy+6YY0sRZ90B8pOgC6xBWMTrmKlBi8dVMJ8
ewyxJ2QiKOJuPwl14D2nd1vapfAc6Hip+ekpF4lkfPHavqlYd1rmP8HfYBqu1yVTzhwXCizhoAoD
kTBuy7dhMPBWrWqrWa+GMC5SrF65hdes94+uk/9lKQXNJP0QFmFJdvvi34Bxu9fv34e64ISea1S0
x+zww+kZFQrngxRIPoiRSNTcxw5JbkE+fcHKdXHHKT1SA1ks1joKm7xt4/Xo2VGBxo3ikQq4k84C
5J+ITtWvoL3T6D7SMZ3HptMDjr+8rK7t/SN1g0lA3lB8hKzMUaVZUcBRLigEdqXsZ9atXgPeCSN1
o2gyebPo5ya7jEg4bcrYSfnS+a+b9OWKbahPMdDpZWTi96njBJNLsxStLceISLc1Kpc11/9Ey6M8
pPK8ABayfVokfaPxEPHWTSHpjEgIF8ebAyQqYE2Nv7r0n5P660skizhAZ3bmV1h1+hUnsOsX3pSA
XKYGIFdp6yNHhdyauwk2mal9kehDlzOZLd9/0ANpjn0qoshJHLEl5E8IoSsvAdR0r3ZlR0TNMqOS
mdNk/aS/dN0dILQ0Ly7qeESlhVycAsuTUPQRI++2VCgsXvSSFdUxPy6oKySCBqj88wBevnW7Otih
X7LAY7BvllLHFEnYcCY/aKKlnCx2RmxLLeC9idLAAdXcFovjAdUYJwfKW9djNeSNqozI/9o0aRkR
s9T++hH/pRiVF0DIFCK3l7i2SFRXarm9WN9d36i5OM4dz9iIy65cFnu7ksNQMzyiChSR9/sN6H17
kNPWk40dEKvyzdXWCgrrVYAoboO2sPiUWCoCfLiItDTnpCINmWuEKjk+ncnB6vcsG795C5SMPvKZ
urQ0lIMZ887nZgEjDmmnwWlHy3XJcIvACPvOn088g0Ok/gtlSWRCsi0XcFm3NIoFoH8Nnp1HpIWe
AtUd82ehIl8fUKTnCAxykxydtrGtbn2uI+q1N1BIj35O7bccf7gKUOHI5sD/tzwcuK3YpdtjWkRS
hYhfeZCtqS7r1mlYNcdBOSiNWVllZ/6ztyBMimUHf3Pik+o07gIX+I5JpeW4J14zCYZ3T2qygcfm
bX7DpVWvjVfKL1cO28PoHSioRNok+4b29o6dJX0sU+FeHA11WZSE8ZbIEc4SzV7ZPzXPiWZxcpjF
f4ysbsha1CukMSNqFuVItfh90wBY/THniKT/N4XYFYBrAK5/P8K/UvMl7MghmniIy/ry0M+Wms48
iFzAvev5+K/qkfKPVwMOOTRYb18pvmbSvqT9N44K1jyTWGBVqhtMX2jT8BEFCayO1iXXA51ACkQ2
X04k8u0a3GtQs6yujijK60x75ahvrg2ISxmiuiQaJAZReZVEA0Ul62SzrpMBddr5J6XCpYdATRwN
JMI/uOaN+mTvQONgB//6q0JaAs1T2ckK3rmKTPYbyRm+PJeiORWZWXrvhdZ5qCy7Yrh2WNJTm5tr
Fxz2SL9d/kdjlQ5S6q0L6GbTPbh0NUrEx+oDzCQtdorobl106Kokj6r4ZsElJWiHlNBWqRcRoy+4
uAbsNiBrbJOdyAcGuVm8atLuV//xZeZhM7ocHqu90PZlGP/reAKGCyF6desFFohrKUJjSEdfMTfo
QgSN5WK6Q+SxGg87VJ3xZEkdGBgyoMEMvuSebL7gjFfJn5XU97GvKSqGfkcDDW6E2BkIjP9QAkVp
volXFYbcl6Xm8hU5ta5AuAXUB9tGlXbAznEF+9tMZINdDZx1o+eXXY6U/BjN3RkvY44N9Xc6G/Ob
EeYs6jgwDyETiq6S7SG/70jBc+TGg7UGhDcQVjEQj3jEGYKS04tCXKOayYpaf8sb5LrD4235X0bM
Pe8uGHb160hHzCbS8FuMr1ahryytgqtpRcfYx4fIVzWpmyQXGtepOu4yOWYZIPMi6kVWz5+pi7XB
PcT7dQvX3CpTyz1G6XNARtX/ctTNQibKq5Zw/qX+tBghxUIDVCflB100qK80BSJnb8W72tR0R+GC
xi4C4M5Z8z240lNd6+eluPlahorGZLMd4uCHvuGf69qIyuZUpphOxzwzw6TPAskGDAj9B2475GoH
O7575Kx3O6BKzHZQ4rS1i5GhNPVG0uqbzlOaDnoCzJooa25Ujmxlh5t/Hxc1kCdrppFKBq2f3vqe
ov0ds3VTr1qi3z5f3g/tV0Mj3fMSJ9cNTZJmII8uInjKXsHuVkiO8KEP+MKn6Yv1PIyZcGqD9r2o
ODggLNOqqokXpob2WcZ6LUsZ7EomOLgX7Gl3lJauTBWNz9zHr3DEBF+vbB0kH2nEdQiVqzFo8dFV
Ol56J7KR2YUDXi6dfPhRYEtqIrUmiRE1TqshCjV4BjOBbNDOQfrArU+9GYUNcSFstEEDGa99VuCt
xiR5YFngrcWjVrHYyOQ1bcrdYWL1fLZwOv7/nYiNsiqwqNFdt1IAuFC8Ug73/foJPOZmutisDnsk
1G7FppgUQ+h3/+HHBVz7rR7yPz/ojpEEji/7nQlmirZh8acM/h7BtY6l7jGLMQ7CPpK0Pnxt9sGw
MvpUvFGzbG1hzY2AUg1HKhIA3bw4b4YZLwGYG2Hzem2htbQuxsP+hKORSKsw3sL5uCuAbMpP4MjJ
vfpmtG/ZUI9jqKjLf4cmy90cUQKu/ecr8Db0GzS7HtcM1Ulm+JVzViWBdK+db9N6zusPhI5w+KmT
1JcpGLC07HMl3QFNg6ExYKVrcD3PRE4pPh9PkTLvFZgOtduG9+qVqV8ca388g/stfr1+JOgVZwiT
MCUT97SA/+LkN5e/TCDslU13XoJvII235GRElxxpPuqG1RtS55pXCKaVu7655QsFJk67TrvFrm42
AmCyFtUcRQ1AGCGyUxOF2Lb8HPRW01GiYgcLl5G8VRER2YkzhrIbfiz2henITnSqa0ezsHOqkCkc
PB7u2U00ByzxkCnk90RSRm32y6ooHJuU6n902PR8ITqnPZyi++FStDCVN52ZsM9QZ1QthHAu6vDn
rSdl+hiSrVGr7T01sXL5gmvKiT0T0VR4fxx4b5X+DD+gqckV1rmTPZ01x8INvLCzWZi/qcE5sQEd
Rktkmi444pTWtUgE2eOkOch9cgLcSxoRoZvVtMQ/eV61Nlo6CPcXRXGdlpdIFWjI00CBH+0dM0lb
DpT4mZMKolbIxKHBdSglMLB0rWvZex3Tar0CBFf7EEvl82tZkdwnq9n9vOIjCxQNOxb67EKVFI5B
Lqy3ayu23eJg5LgSNROa4PZXX5AkG5AB/SgO077KXWdj/unfomV59M6lNhETeyuz97+diNQyTeUT
yxYQs6hscl6D/8ymZszclCLuf0RWrLJ+bSqlBKSXi1HkDV7fUwux1U8OKoKnIxWfRLQR2CbiL6Ev
qQ1gGnoB2hMlaeFz8KTWoD3co2WvUdiBavJhvy6gtqMX+EbGdeztVw9d4HeVqTlzJLiIFAUMPGKx
qoC5o0RSufrBCqwlXGASqsA4Bq4A+CUFDA0u3AJfZmMHUW2d6VEjRXMmhMoALWboRARnhv/HX1TW
c9NExgymx44/Ba2rNw1SDIOtIqgP0Kp2CD84mDoFvH0t9P7W0/vEJ3Qm/m1oGsRZ5nAS+haozwV0
1xrYWoFkWcKm8xDlDcovSM8m6s4OU8xpQT6rwl2AIXTakzhpq2v9aV7Cs5No51tAB7nDO/+lOiea
Qy8O6rAkw+WoYlv4ow2yhDyde6Ufd+oCVbzPB7B2VcsoPfX0tpMRJqANu57Jv+f9l2Ro74exGXw/
adpZwNxHE9/Qe2jIAGp8IbCQkSoG2O/2BHD14SDvwXkttq6FGoxgPg4QCofKG7P1DK2jkyrfmh+M
JL4+SUSxiuVEBZ8=
`protect end_protected
