`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dToJHbXRVRv96E5wPK979IW7dfp8EjLm+Juf/IVEmFkFjuiVQqQ556kKiwekXKHtR2ViKlVIkHpk
fSrr/nO0yA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZyXF2JLzD9q8YOAegjTfR8RM9ueUqZW5UqgiOPFe0ZI5WgheqH7grm+BHmjq0raodjwAoSWcuANa
OkvNOq/Y/Gswq8qP9iez6WpVNY637d5szL2u7PUS7gz1l45Ipx4BQe0vXnXioZoykyp1wplQdhD1
u0/Z+33fEBdGp4e9RC8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gr/LBXTOczMIsXMjsldIxwJmZSpIdz2QZImc0d/HAMT+n6QJ3O5xY2He5TIDab2seuCYdn7LY0gq
oONrmkdVeuhdId+nE8TL1lQ2wKZMRhXStSVnkYFMNpq8qoqCVyAvBqY8qojQvUSYT/yVJajZM7ya
c9anokkyWLzXZOVUh+8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1xfQZW0RyoKNOMWHqq7GA5MYDWJNFs/D6C0MBpzo8LLW/lex44dODJWpsiXjnKO1BnDxdIzZSuMb
magQML+itv/iUcsEpAhgZ4SnshFdKhBplvBDt9Wrrq4uayMiExeFQjb+IZR2IURKYCbH2PXPz26O
bs/5dX4UbTN6+DB/ph3Vkju6KfsiAW5t82d1mMJZCYazsvSSMYF4Qsj2/0G+d3zS6S+9rIQGVc/k
DAgxKv+56LmUTiqcL2PVAC4Oj6JHw9fxvMegivn13Jm8eD594EBeb7q9fsrmrI+uAHcGr/S80yod
srIn5OqPYy67EMU9XpJnyYC6TBG4AdmK0YtzKg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dDTy8Tavz5r5AdTl2WpseX0f2dL/1rIAq9ekTFPNermaoKF9kHdYsTfk3lSEKAbMOkTkbFo3Rv8f
jP3jDvJ0MefMulnZPsm1hV11ZzkjxXLZLjg+fLzYXmft+FIm7xJYMwdjK2pMeivMUuRnP3KgmDOd
i2GOh0+nwJJhI+zDgkJc/uHou7HOi7aKFao9YjJLmhQKMFmCoqaOdJ9pco+VWzxAk6Mp3hkV6JWJ
dNMUEaeBVYRfOYZJeZFQKyTFBYnGd23oZKccqqmRJhihzgbKJNtmtdE0NVYTK2g0nwBHRnPE0BSp
2wEH13eBNJkE+UwBXRAuZscwkpHgPfwETsbeAQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lRcCNvUUAu59c1L7bFLzwafJ6MoNu9qZgbX7ts4JGrLdpyYrwN2NMdbi/Zs53UD0oS7Uxy07S+Yf
TlQsusSfzJDsy4FrMmv9+4oGcbVkhLOB6M2uK/YBOIGln8ViM/kd3muEKt2jw05Rkg4zXEzqSqId
+jqgdBHcBsEgiGUQMi/Ir0xZdqXICjKNPIX5xL7jN7crHvy99DEy5qlt+dMr4ulhQCW5Afcw5d1A
N6wJ946Xhw8qr5pWMS2ZynobhZ/o0+5wtUtV8xL+C3Z60N9fQ2GkQQg4JQTZQ/4kuQdEMkZcj/7f
ge19udWKONXuiWbmYRQQrNEyJzylWDkb1tIeQA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8928)
`protect data_block
sGK4JTBNTSxebPWFFtkkNqVg3RG0GV0eeGDov04vSkVVKpy3NLyQgGljTZkxGaCqX42CyQhUdvEs
x2eUQF41hxIbBqLdV8MQheaEpSC5nWDE+/XxRtTo0z11lCVsbTIBZmKBN1+HBQLYL1VKuR0l4AHP
UCoZ42JYZ5Y4bTgwn3Q9YkS0DX7N9tFZHiePkEs/HH/Xu1U+XId8KopHtab1p6iB6Tv3OEhc19Kq
5Z6VMz5xMBRViA9Epz8dugtHGEGpyuvcrWnphOZ5Lkg8E4C9OtlnhJtl1vdQ5hphME0EQlOZSsR3
Y53hamnAVIj2ZZlNi0za2RlotJLGtRjPOwmKfhsasleCyQMSwnR8FTelU9K8PDQhH1+qEQCKXnrI
3Pxgc3TgvkdiYbgKI2EX4ZspLx1W+QEyfhrikmcfTd0yhSVeHQwSpyI9TqaJ2g/YdqkXj1N1/evY
cHo+8CSLPTPH6KlXJdIRzIZzRCG28MFEzyZpyGqSrKjJa7fLViLv/Ld7DG0TJAHtMrZH6OKYTD1J
X+jQO4WtkSiKnGcbuuYcWeRA9dNG25AbDdvguBR/XidfoqsJSuZ859QsfUX3f93X2tKOB62JjDHt
uKakGsxdl9JXADnt9MnKN3MHslCIRjAMZref9NB+cmNaB4Av+zjHnEFrmi4TDW4+acpKsFCjPnIr
wDxclnpx5kkzSQVCOFKLe0kGElzjGuL/L73i4hQEmKs+Xhw9BjBik4nhH61a6gRtAvc8Ng0ImM4P
lHjd2xep/3al61ICYElkbaLXoltgZ1/YbbcUwOxUBBca/Tp0kwISd9CMHtARICnHFrQImXRVacLg
giyCp1oqVEq9Q7qhAQFEsW++GCPgQocIxkve9YfwkFTjFEYH2Vv7QZaHIDkXQLj4iVvCUt6ZnIfW
RJ9KVa2+4mF0QuT7qX/MlEC77okVNM5AivwNxRw8ZoKrMM6CCZuhge91dExglbQzHjEtnM0Wyl2K
LPWvyPwe7AsXLUOhD0C1PV9tqHCf3KUiCKtNi5ClPDU2RIlaag14QNjiMcceb/lKuMgNC3Q1yNF7
HFzpvV72GLvHqil8NYejYuw4VXaQnZvQ/jd35oETZ1i7qOvC5qy5uWtWi+56W2s4FtcDpUAeU7ZN
eukIgLL+7VN42U4smhGi6wivtob7U9eV4G6Tj3w1xxuc2xqe8Sjt/6N65yU0RQmCOdNBkHuj6FjR
St0AWmvV1hzsnBLZktXOz4xlO1rJ/8i73o38YaGWNiXl2UtvP6bwYXbqdGifO+HqxXEa0IZepw/r
RiHP8GervyPbgtjEQXFrKagBvR3NjiWF8k2cKv5jsN1Ew/T5nq7TfdCh9X/isGmmzkvuGxetJGZ7
AKTba9g0skWt31ptg8xaZU5YKZ7Hlh8MBOrncO53iqD8u0uPFCS+zeLF7TPq5g+Jn4BAXyGgJXXv
AZr1XKGSMNjQnG5nbz6dOGsqzAnFG7meGwuAJz7vV2kr7yymI8BMS+v6+3GJV6B+HycgWnQ7MEfI
y6KBDb1OOOrG6c2WNw8KvlUSvVPhtZKgeApL3JoBFW4T0UMp57xYqZMja61ym8rsuILLrI88SQGV
L06oZHUfbGGNhO4NCYmZwJPmVPQ5t6N6C7ReBwfKRij3Pn0lJIHdEfXLcIx/i7fd3MiE8vSxwc4B
tbHBNBxKcC7Zo/inGG51SSYhZDuJJgfEEUv8Cu8EgFCkgKS1cBBQXrFMklO8A2oAmNHXwOcZGsr/
UJ7DrmQjE3gOYxlRc64j4nR22hU4Dv9PF2fKlQ3GpEGVLix8+Mkpv6p794ZHv6Hv8HNN4opmn16r
jA+55j10IhuhgBb40mebIhKkIbss3jbBodkrI7ATYKvLJ06X7P9hE2yCF3fZYGKWgix9GZiSFG69
7S/xF4/ZKuUt27dYGhXRi35ecfeIoxpbyziiR0HkoG6n8SlBnDCr/1uf1Xc5TUjj3tcaQSThQ3qv
3nQ0pfTsfvR2gdWjxM95kLgZ2Zhr0Kw/w0WW8ZHEGoAuxzGv7byxOKy8r6aDJuzB7VmnOeYA4uol
T9PR6oiDA0YReQgjG/Me/kB1j1UsDmnT2taNrBOsBS/yWbZKWL4K/Q2sx03xpYMbHpoRTTS8jqCO
rLx/A1nmFLD7zk3jjFNLBFwRJPLF3neTDcmYhoPUmbnTkqb19JSXZeegBAs/RfTkfH3HgRi0HOJN
JSY8HIQaS2qXnPnKzx8/ExEpZrpDPEBH396tdsa0wledfrEHMsKuff8RTSUlDLwAKlpo8lJts7uH
gt3P7oyYYUYsmetlavVOkJpCFc001r2mUcB763jP+vJ3NnCIwA5CNXxGx3MTBnGRA+9jmH3QJUzX
iizPjCWpsCKLvgVeQGrJuhIH/UV/vARfK3WxDx8Jn87ios4A8QBzWFA6oO3Y19rJ4FMm+/IueTlt
jTJiAKau46D/lrDNKUThrJx9MHYlZ7kP/C/zKRrM2/v+kEb2zkKsT6ym6WR69mHdRCdKNoBNMGga
V1lOun1lJM0UyOr72p1ocgq2Q+s1Ie/aWQnNtgOsALUWBrusI9LnH5VIgMp4BtFiL8ZiAHIcEL9+
149AdAGarmtVqenDC9s7FX7/d3+PS/FCd2A4eOH1+EHEa9xJhvmafrUVL9SdewsrPEmMnssnTYIP
x+nghnYoLzvyxNGBlwceituEjXR4TSe4KUhKBZvwZBT3gMqqG57rY9qsju7XmxTHokoOc+z//qUu
gi/d8nY9zqKHJK5CAaaOjiTaCsXxD30P8GZJipXV8K/NQv2QeZPgCPU/PtnSyvX9ATZ7373mBmSW
4bTaaPMqBb+MeR3bLowu84bzr+OL6QXZXmboDt1VZQOq2Vd5mS+ZI5ckUJsTtCDVqV/X2YPvX0Tc
pJ89G8TUCR7yVTt7mmPEvKnuOGV5KInGxkyTD/q8onFaPkPgENMtTgsuOlZDDRnhOBRvTGmEvDkR
SpkxEgt6A4UL5msTFPd739+CH2DbEAsoMJnKZ7WMINVAlVtgPf/F2QEB0Rd6K9uFJXwMdgxwkn4t
c+bDHclrH/81Lx7RmPEQBurhSn+p+aqyjKoMcLa/rLxoo1P85lNyk1bmE+8Bgg2xfKau1TWL/cyA
FWk/qzuY04jDcwYhEYVrOVCzl1vXoLvF5KXn/FpaRga+z4+oF348ZxHgGPpuoTT/gsFsLJfj2NT2
zX15rzXNsNBaQEMB2S80WI7YYw0trsnbugEXCs5O6WKe2UlFm8a9v265MB4hzN5Qf3HVP/rI8kOt
xMMCs3uO4ilyRZsEMUrK+r8bits1Ezj9kHRI5d1PbvoU8d81uk55CFnOesuP77+A5/vqt7XGY7D4
tjzQ6cxDZEFmVLHQYdkQeirDwqh0kPZhtMe9KHbi9YPqWqX5BYrzSGhKqzWhzI+iCI/F0ObBOY6A
DNiUOb0TvoZvYhvZeqzNod0ym5cl5jwtckh44mWDYqVjoGgZaxd2F/vArJOCA3B4Fgs/8QUPRVxU
6gBAbalYqqhGH3IiVbaIsClwl9V49DDY1cz2LmX+7c+X0YIeHE/NKuZQdRQdkZuCQ7G4/CSkABOy
LsmeoXhyizwu+fPFl5ytSHcLZN8ZB3LbS8eFuFwZ8Rbwg/j7zjz1YCrZ1RIsm7TagEjH4kGuZGm+
rTh1tRTDjgigvyjsG5JdhAYwFdGiHrzowgiSvzHEuRqqxqNGy+UvkMxDZhA+4ew2pAYsMb1TM5Mx
zU1qe2hr3+F+noaO6YQ0Fux1I2lJNG7Dr12oWqjjIw88zBzhy7ka8K42NVVPa8kzWnepSs20Hu2/
tQlKkW2Kt8fg4sf0qUAqK452G3CkjvI8X6CnPScqyExgyuBysTbcBdHJzC3tCOePXxGxUZJxb10f
rG2gj/UwEWDVfDzfKuC+xg15cbKK0o89uiIGJ4hHB7+OQEPYZT4YWB+pDBqjZtUbzbmnvnBneI9C
g5ltFvZ8/e9V8fKaP0cx/4ZxzJIrJdvKVo71fyaoUA1zJAOgfSiJTIcm7yJo+tlSRB7sD7XD6uJR
9lMxCLK3uBKAbpLqt/eH55D521r1luKot59jzTSLUMrLPhnfLeEP25QVOk2MfVP8cPC+6Cjwlalm
XvU5owydAaR6Oyc4hHitKBmOMAILIj+KgXfPhGdpLXiWKyZATwpretf4BR1mQYJrCT5a+1YOohSv
xPw89LuDPQ4IoStM2fsLj68U7tEOscLx4aGDGnc4mC5qlaokBpXyFxWbeY0c7K50/0aZ37Egb9ej
LQ81X/duCxrIAqXlBE2pn9gUWz1aCyyd5V3Jo+NYuLDtJsy2oGX+ajEvLyZxATPna3JnSFy7JvP+
NePC95eX9jvpeQLsKoYZWifBbkTg4Vu9RMpobfKHnlstMOPEHLMfB1w19zHKC0oovKLelGs2182u
sfKwJAHgpB8/E5MmvjitgmIU75J6f8AhWEx4D7jnbzoc/UdsMmvgn2CT3Ldbq4ZYm4YSx2pm80Pr
gd04N6lm1NR/WduKShlEIOXoDMJl/6bDR4RmJSsrMnEOqZT7gNotS5Cwvg3iOzeyl8qhIvYZNZeR
cJ3IrtT/hGmpXpf3RJLnHFmAAhMUYQcWFpedK1ESTlmNTSNo7I1alCjQ49IFjpWG8WebNl6InSQE
NOzTqjpqFYDHk2dZ8ILnTbJCr1U4m2EV0A3gdgkPrFVqvhNv3ZlLB6360KMQAVymElz8iEGJ9n94
BZEn4B6/B0UYKOIlT6fVNg3kjQasBygSsz8iiixjxOnWkgwm2/uGWduX81xsLe1hga7iQN0vvc4B
8Z3lpmUQlRBGNu5egMYNTaqHquVas4yxiVQcB+uE/+z5TBQ7yw1GnHQxzHhC0mVVQqVadwpUbW1i
fOgNS0Rn0Pg/a0QjsHV03ezR074ukSILZxPy8P4mRjHvqG21Eaj+TXSkuymMLS8lQJPqtVFn0nhK
EMrq+RZyvmZ0ywwVV5EGQiLxz1GTFmd3Vt6ESttG8bjNYdMjg4GfDlNg8R27lc2V4TrlYk6J95pc
WWx+kZ1Q/MQJ7r+n8znhuyYd/39TYOBo1Dgws0WV7vxiiIyRMP0sIXlNQuYlZmMYs6hukMpsY4T/
FTeMmW8Oc6OAC6QM2mR2OnnbKWW12Jm4MHFsBp2MSPO5+rddBnITD5N+xX7ULIrkGWd2sbyIvqlV
ukY1rhBpoWqkFGJxhG3otTh9TUmMaXszkIrW+gbLFYKgcoTRVK8thg1PJrmZ7Zehlk2ruzcyvccw
JW2BpHaidXahS7K7kmxvzPIJQt9GNs1fzkVnWQJEbYgV+Fa20kIQhpYZF5jy7hJZj/9apMisSGPI
xXOev9hUqoOCZX07z8Ei/aWsiRtE3wRfGLbcXsOY7paxvLxo8oisbjBGGqKCdYBZwwanMHEfM7O7
j7vAswDAbQndtSs1fvMp9q+Htc1Xzxqtr1OQnO9gOWkS04tM7jQMgJmhoKfPCFYA5QWIC0bhfmEw
9RflBVahBKcbK2vsnQ8O0yFDsFxVhBZqKrLs8c4yHePyl4Rgybw7C8keOUe3Kit2p9owLv291LCw
MP7ulGufH9HU7hDMRDNAt7kLeIUzrsJmk7B6zFhIEJQqyJ1ySdaQfAdvhiVtrx9sDsysq5u0cb2k
FOqLdy1qNoMqm5ux28DK5+r9YYpk6n1Bmw80fKPLbOrT59GfYiACQrMXlBWJ7Z/lsHg6vy37vOwS
nqRySdAmbV7KQcybuAGnpcjomSBe51PVyxXq4zXNcjw58BDcd2yOIzAPzNTGWsmxgGYzXWycLYtR
BPukXpHdFwTiKU/8HuQaWsjSVjNNfge8UvSvfOn/3X5p329I6st8yj4dUGkalMA6Ivi98y5p7vuy
eMk+FPTrUTHOCqph8A72CdgnUsgW+UJCrNa6rvuSvk1ueclTzy3ZXyE85/ZTDbwvPVQUN4aMSjbP
jMXF8HPuVxNGHKHc1yljAPiEfRIouqA9WO2HE5SAmPXbA/U+jUC5JYA3OJlertXGzdaRfBjlqOzb
Mt5P2wT5tf45cBvjW8jdzwypLEkRC7mQChT2NFVEliYrbz5/4ANKAPjhVh4eiOefLgRsVDX7XVCv
Z7NNlX+cD3i63HK1tEo9eydApr0lpO1NWKtHIQxW6GXveSvVZjlSCAb/N3a3GQEjNIeG8VkcdV5a
1GbU5HIQI2Zpg/XusYyrlMufzOrkh6UKcIsNmDobLwgQkiCBZ5sQOfZiZHUrumqR+VVa+Z5lhE3B
aDt5F97FM9vtpCYrkmEaDu8LT7ByZ8yYD06pHAeTtFGFK+yNFqMHKJl+U8y8azEU32TSyPU18Z0b
Z3zJ6PvGEN15Busnrd4C7vWUrg2+3yH1C3MNjryJrODaKWVHuJFbS+E/cfMryyqZD5ON+UT9bXTU
/UGLEbICbM5dSHrEMGK+ytX5RjGpSuPoejpZEfJOfIzdhgDLvBIzyJWhqVT4gXXSHlTkR5CuN9bt
Y1vND3H2uVTEaTtqWIp9BCa4vT0kbv6xkdMk1EqkOkRvCvxTCla8lDJNf/OlkSNt9IYu1yJLMvFx
/W5q8VMxubufxXAoMFKbvTx8T0qloat+mg3p94h/vxRSk5LornM8ViAL+0Pr7nXiLSvI1Cb8bVbw
3QyjrrLtOnz4aI9k/+1HwPDLUbjD4wBYtHynp0hgS6hozLWSoDpYnbsErgoOIoNiKz4l1+j00GYq
kkbOvYFfXtynW24fvbb4+mxcdfRvqyvLRVITs8PLSiwxC98rP5WdYvvwQNBXxljDb0brdB1ZuIsz
pwjvrWO1rRuOqoMYgr4jYYn+/ssslbOtqt+nz1FlYbiOOiHJ5/GPjRgNjcekIf5HlJlcSO9fy0ud
czH/GkMSC6axLTAa3MxQDtuYdJIXvms5VgXTZ/vmcZkEkRL879SHnDXwtJ0m6wPGww3k+lvl8LXx
Pgl2Mcx+ADKNJqC/EehfXRIB6pfbsBG9kgrMuPMFKcRkagvqlx+spOdKhhRxpkOt0EX5fwiJ/Tiy
EF9UGEkUruaHoWsVxBfWrix3R4ADc8INTsQvO8RXK+pZgeK39GTDOqB3HxIMmTnG9saGmnizcrPY
2O7pT0maHXaCcmJkNeLTniN7TTtx3YYhWIKMRDlikD9XMsg66eqnQu4pcsR8MK5VpG9Jrp7ppknY
Nq1mmZA38ZGd4RAFxUS2yDF+mVDO/Dr/u0m54YSXvv8KiXzSwnGks00pSy+KjMbvF/0jEBEjERaX
CS1UVvQjLTEiMEBvOFLwJ9l+0Qy4i6nu1ba+HUbXU5MiwF826JImvBIa8Q4oF19SQ61272rTwq2X
ESpHyMMyydzv18yiXbl8K7ACwJKszgCTHEyP1EqqtbGmJWwIIXtFx8jjyM4edNM8/M7NsbsRPZng
F5DzPnabcl+1nAZxiDjlo+d5yk5ZeazfjDMeke/f7s9oiuT/S83LddMadD5Y0mIDEj5QcwpKij1r
n4BCfciOdEPmKnr261h4fiQJon0JHybyA09WkKkplAzTzzzdRD7VaKJJrlgQG2W6mkl8qdSLwkTe
sKYYEr+dgXkSkduCHhAiv0BN3eWJ7jd9hoZdfUD9FDUerMAogv+llTxr7mCCSK9uLkfPvB+migI9
01hYnRU3kteNs0lBCQras+bB5dnro12hFV0mUc8iFBMoEckiHwJuHzAFctyxv8JLlaxhxLmAWMjJ
ALcoztUvtUjlOtEYNMzJghwO9oymB3IBVyV6k5UDUvUNOX5i5DRQCLHN73a/Ch9P4GG/fQ9wBpI8
WhyZqmegwrXnTpv4PkJ8UDoN0OaCZ4x4g6UsyaHgyHkUcsdzTv4j7hC0hkBhuGX0TxXaCCFfTiDh
/szmK0dTuDXRtuti+bDrCWxeRCqm5yGtzuXB5pnc80XX/j3EhlZgJ5DD8y1aaF6IEpUC5m4HEvjh
jEsm8FJPD5GuJo+fbBMXu9RS2EnRBQxjDrszfxyhnaNq7OJc2jhF6ZJBJf/GqtAatxF4qSnpC9rU
KKAYJfmhG/ufhn4uoWHwK20FY9sIKDs9e95LBGO+4BIgPwqeZzNK678XRW9+56leD8va+y9flvq6
1Emetlo/P/8oiKqatnB0LsGOwsoJaxhjGA+EZfBA94aEbs3ui1L+JzfRKBOWEBozXtmrBWS9KhKm
kdMIdlWNGoEQaBfIQBcedvUTSUzEjs7+5wmnGoRPfXRIMVmrOkYrW8qzLzm+lUvPE0fa6SvLmBcF
tVliG5MDNCjSOQQluiQvbIPql9B0/XQZEjLeXkhhuVFqxSSZ+Su02XBRjOy3PFyqF/A+gZsGHpRA
h8qnaXRSfRcLiz8jRvC1Q9ebpor6sb1n+f1Ncv+deImH8fIohaL2LS75QZ+1v0haOSKkg/s9D76w
VOC9MbFc+Ebd9Je4iZFU5kmatqe0MF8VOQnSRI+kKkpdaOpfAh8+D0AfxjMDCjw2bbAMv7udo8/i
0k1VCI+V17Fxc0rgfMo5H1eWm8DfyhcB0EQ3/7YjhA9tUSoj5oz94MVZoe4VGMdjGOJlXUnAUcg3
nH5cDgUvSEYCsrkiAmbU6yYV7hPfrMGWXquJh0cVQyLtC4kpEEQ4+XABqGAth/GhywOTiZN0ojGv
GUPS/WFLbPE9xb7hd8wJxRnK2mT5Te9C4Wsyrmu5o7St9Me+DXPcvYr/ZrbWOI6dJdMkr+QP+aan
95JssH1SwEUV33tytlkd1cE4SLGdtWMM/PDHyYV7h4HTBZspUGEfIRFquHpW+wlu9+K2/WgWrtGx
a5EyRCRKXZot288kGIceVUn/BcDvrFVY1vXlcom5nLjfqLDxsYwDUdIZkE+MM/An0w9GEg/N79LY
R+fgyJ+mEh5ibQw5mV0a0hjof72HzR74lKKYHa46njBB3auMpgv96nPA8Yrdnkk1+yuGjhFR7fJw
iQY+WUDF0hjsTYCyyjNtrjt4AgFIFWfFb5peswOqiWhqDvAw2of9xVG8LZ/c5zHTEuzytNiCHeZk
N6P9aT5mo10j7OH2i74TVCxwiNKur8Zd0dipxCknCSiotzGXP8QBDqffkzuKsbQFOJzbn/y6XH03
qREJS72uFflczqFjZ3gG1lS3gnpskcGYIbTn76rUI+Q/Ylb8VdbaF0WjtEn7Pz3Ek4mzIQRuPuMt
K3+ptUNm8Y2Z9pFFHoMD4DxL+k3DDt0rOabUP70iPEvLg2MjkIJutXlK0fxFahPfEgxBsjO34hiq
NR1piYM3f7DwxJ209YMxqMQcoQVtLteLov2XuKlDDshpKSBFtoMYM4voZcQog2wBjGa3/UKg/TuK
7Cu8p3B6j5b9js6ohQBnxZUPrYpzKgUaN4BSOnjS/WEZKSc+XO9lTrZtdR9steRpaWNGR7/+8rZF
8kzSsjqQCype1cfsC2ojAa6bRIG8CYiZ+mv5yk0fyofLKKRUkolFZr2boQPtENXobY52GzHmiQsT
WeGYvDY5SVrm7cKy+Pycd7vmKt2uB9LibaKQTsu6uTE3DojqC4Xo22y0pvRzH8F8IEOcgmMpigST
+oHvdBxN/Ef5mGdE3mGL8ov0a9Bvyp1CikywI4CptxVmtMmHwuJ4BZi+WW/hvAue711HVEzsL5Z4
aoVPd1oPedQIXcjeTbSgKpmuVl6XMamToBGuWmWX0wWN5AOBgrEBZEhZ39eFe4U6NEVGD2URSX4l
t7HQJBA5LALUumgPNRBVQVjs2lPt8xDMGjvK3Z4CcrULgjpJvGn9MeXjehw4R18Bv7hoYQsSic65
pcMrv64JEgYUY4Hf9n/phZToCRKupbsFkXbDvnTbeLma6Qyu6S0ESC59WUTpzcnzST6qzJbjMTI6
PJ1/Z7Rewf1Kl8+gZmh4tpxqzmi6kgXByHkBOsofor4u+sP+ssAmdm9P1l39hh0PqS6deXqdNr7X
m6x8Mk/bM6EVtbYFw+q2/ZxuQc1G4icUNCw26WEdGtLNYYKJC64OeqOwfdij+D6VwM3bL2izNEoP
xLpIq2cPHjDk0bEFWVroG9GMW6jUmDVLisQ6oBgVPxMzXPFVtBH8M7SRr91hdonujNgM5LGlMuyN
QbueQHSseZsHdI/Kl/Jv6TpJu3Ajln6dMnBiMGXR5t4cg4mscpBjohz3g/1uK4Sct//AsEUpt922
lu+fcNAqmv7G0MolL7bXBf3djEm5J0dtZ/gagQaLRZpvSJw3vsmSmthyNGnu4rTA7SHSeNI5/iOY
B807ekxLAqUAzAGOYfzgiUC9nkBZ72uPozXvV0dVtkb8+cncPwrjW31E8m4Q/EkkhG3lbEUsPXMR
/jmAVmy+DE9vEbw+88Brh63t2YIjAi12PKLg9uhYJvGE6d0Ximr4iBUWPFotEYS5eFgrUwZ+jeUD
8dSYfnlINi/qP+O6qHbqMnHOMdAYZX3RhL2N2YHwa6VzqAIo5/qKJyZTN2KlIK/Hz2Brhx07Co1r
Zz1/ZcsDXkt8hvnwTfrtcru/U4t/js0BoXALLnemslzntRDS8X4W+sDJDMws3doU0UmHs9j8TtYI
ToBYqAufIpV+nACqpHwYa742FopxN5bAxy37I0YGuZP6HMTpYCnCLQ75LGRPdDV8n7h5pzn0rBu7
+OoZedcwovBsmlwzNEV/Du41yshyYcpjJPHNcov6E7Bl9DUjCkanxMUmbfbzKNk5uE7wEqeI9rVU
wCBcTGBLut7o9fB9VQiMoPhKgNz5FTOjD4+Iba8OAmXmZq0yhEqe0DhiLzdLFUukrTA3iEMfKdtD
hChiTWeDWR6P8GtMHSJDKtseetHABzJj5LRid8VmsIv2ZoO51yaSADJmCjT5JBlzZ3w+Sfbdgir+
4vFEGQtJAAO6dvaBimiXv8byRZ13A17iBYkihhgrssY9ejtVWjITtoUHDFP8e/V0CiNXTYW6KP6h
Bd8vv50hFjt6OWSRLKt+UgrnqsfOrS3kWTkD2QTV3/uzWCuw4VmYK/bR6GTH9xVG37ykTW488/AO
OxR1VvZgFgOQ5BLujHOGpiVumFHeJ+igOWgQGQeBnZCitP0Y3LE2PAquoV1a9y1CclToL8q7WMyc
/VorcteG9ODGtT9N5nkkjVV83zpSaSnDcxSRGrYOGWtEdWpAZ44XXyBrXeWmny6Qf5/vDJC6Sa3z
ZrYVR5w2qQaNeZsOQ1eTHmvbNHvbKoBaL1UpNtuUHvf1reMcqmDD7NzHUQg8XSv2mmafH2caOfhK
CypoRCUfcAP5nLzQXCjreu81eRm6G8KKKyIVUROz1LpHfz/KIwwSXrRYdOeXhvCpbsrEsG17hRsv
ic3b/UX80VooiCldz+Lgdp4BJnz1sQo1dOfy6cVaP/HFikt4DLLWsUk4zZBA7zdkXqOzOEcJh61g
fDCo7nT9np1wMGyvyHh5J6RdQDQeD0LwD5jDdy6HH5LgQoWZOjdbLTSxekx/+v88Akn7gcFQSbHl
Eb0xr6d9pJYitPPnc9T5vJtStpGigNgORmqFsA1Ttr8wEWUOvqLSVU19JzqALnt2UKv6MCr3R6WS
TJfbQ/dMCGJDpuK5bCp5ykukkeRdIdBbol2bQb0385WhTpy432xuF87qACdGXx8nw/IHmpwX7Yjl
QMzPLKrX4nhROgeKBDX5hkGtJw1QTL6m1tsyCikwAL5VQMeQCelIB6nH7Z1aX2k9UlFnVmo+ZaWm
0SStaLZGQ4bzQP6NnFVczJi9J+c9K5+cOmStewUKo1LUmVHwtjcY/yjoXPRJw8Z19QrtokwaFMdo
3ElBd2trqxLfCCGIoxURc/kFPAjuHPOq2v10ptA22GfGrCRD34bZ8CaZqkWWs5goKqrcCfLJouBL
uxeNlX38npxYI6wwXhKGFNxqtpMOTBjFjtCBoWMnC7p+sWwMa0SPe3tOdFmGzArAWS9q1yZhDHNq
+r6HXl3ezDijhygnUoscjEEuMIHBSM0kl1LK52Cl3l1RHlBO
`protect end_protected
