`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dToJHbXRVRv96E5wPK979IW7dfp8EjLm+Juf/IVEmFkFjuiVQqQ556kKiwekXKHtR2ViKlVIkHpk
fSrr/nO0yA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZyXF2JLzD9q8YOAegjTfR8RM9ueUqZW5UqgiOPFe0ZI5WgheqH7grm+BHmjq0raodjwAoSWcuANa
OkvNOq/Y/Gswq8qP9iez6WpVNY637d5szL2u7PUS7gz1l45Ipx4BQe0vXnXioZoykyp1wplQdhD1
u0/Z+33fEBdGp4e9RC8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gr/LBXTOczMIsXMjsldIxwJmZSpIdz2QZImc0d/HAMT+n6QJ3O5xY2He5TIDab2seuCYdn7LY0gq
oONrmkdVeuhdId+nE8TL1lQ2wKZMRhXStSVnkYFMNpq8qoqCVyAvBqY8qojQvUSYT/yVJajZM7ya
c9anokkyWLzXZOVUh+8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1xfQZW0RyoKNOMWHqq7GA5MYDWJNFs/D6C0MBpzo8LLW/lex44dODJWpsiXjnKO1BnDxdIzZSuMb
magQML+itv/iUcsEpAhgZ4SnshFdKhBplvBDt9Wrrq4uayMiExeFQjb+IZR2IURKYCbH2PXPz26O
bs/5dX4UbTN6+DB/ph3Vkju6KfsiAW5t82d1mMJZCYazsvSSMYF4Qsj2/0G+d3zS6S+9rIQGVc/k
DAgxKv+56LmUTiqcL2PVAC4Oj6JHw9fxvMegivn13Jm8eD594EBeb7q9fsrmrI+uAHcGr/S80yod
srIn5OqPYy67EMU9XpJnyYC6TBG4AdmK0YtzKg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dDTy8Tavz5r5AdTl2WpseX0f2dL/1rIAq9ekTFPNermaoKF9kHdYsTfk3lSEKAbMOkTkbFo3Rv8f
jP3jDvJ0MefMulnZPsm1hV11ZzkjxXLZLjg+fLzYXmft+FIm7xJYMwdjK2pMeivMUuRnP3KgmDOd
i2GOh0+nwJJhI+zDgkJc/uHou7HOi7aKFao9YjJLmhQKMFmCoqaOdJ9pco+VWzxAk6Mp3hkV6JWJ
dNMUEaeBVYRfOYZJeZFQKyTFBYnGd23oZKccqqmRJhihzgbKJNtmtdE0NVYTK2g0nwBHRnPE0BSp
2wEH13eBNJkE+UwBXRAuZscwkpHgPfwETsbeAQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lRcCNvUUAu59c1L7bFLzwafJ6MoNu9qZgbX7ts4JGrLdpyYrwN2NMdbi/Zs53UD0oS7Uxy07S+Yf
TlQsusSfzJDsy4FrMmv9+4oGcbVkhLOB6M2uK/YBOIGln8ViM/kd3muEKt2jw05Rkg4zXEzqSqId
+jqgdBHcBsEgiGUQMi/Ir0xZdqXICjKNPIX5xL7jN7crHvy99DEy5qlt+dMr4ulhQCW5Afcw5d1A
N6wJ946Xhw8qr5pWMS2ZynobhZ/o0+5wtUtV8xL+C3Z60N9fQ2GkQQg4JQTZQ/4kuQdEMkZcj/7f
ge19udWKONXuiWbmYRQQrNEyJzylWDkb1tIeQA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 556896)
`protect data_block
sGK4JTBNTSxebPWFFtkkNlMVovOua6GMyIdLpjKZx5Kr0GFvMv/+HU60T1AkWZxsZC22sQn+X9rV
T4qoP6Lxa7Gtm9RI4TRaaaowDPPvcLuJ9B1p+J8SqyK3Z5gUSFWnrj5xD7MnkuiOoLRwZzElxnPn
LS0oEeY9zIimWUwDVNt8y55lTMlgaqhGT+KAOjlDv/868FrpEtx0e+j1+xAGPqieFfK76XVrGpnn
irh0ScItreIvW5ubuNXSCiECaYs/vy0v275eUwh5elDIuCOc4b7sUaeandzq3PqcOj4gErfrDp10
7I+rcTCVr5TiZWb+HELtXabhKCv2wv0HjIE7hTYgJLNrJ0W9iwXCr1W52fv8b2AJDyce5S49eYaR
wg+sih0hXyJely5jPPnFI5QUtvduB1haYIN28vzBBn2gQv2HxqDgAHsdhK1wDvvNZ4jx8X/7qQbY
oHyGywH8wa4UoIu9Qm08lSzsN+miGQNBXdR3X2Txac+utybx7XdO82SF8yIPvZIb46B/1mzwUukf
en0iXwqNMJDMm4r6kD5pjawE8mqQWn53ENp+4CWPehrOryOjY26YpEjiRTXqihEE4HqonFLUbdgS
HHjapKI1zJvjLp+lKw7+cjxzCwC3NSTQQPUdKRlUMW2bkr2hpyWNftjOg2bRBtLTilS5+4lkecj5
nVdXY8u8f0wCzycb8q6v2s0eK9esqcactIAuWfpsiChUrvyCJh/BaSSoZg+ttEpTiXwRdF2bCf0d
W695N+08TLhTelBCdQdP9jBKIDQVbBy84+C+7F8vY5kEZ0roxmrqftdNpPhoZaB7JO8K5Xc9mxAn
v4ChY7DLmzDcmZe+b1D9q56XtBeN6G6tck+KKGV4A80+5z1+AEDGHH4bjCDepRKjs69dNGTsThHp
j4l5uJDj7QnGpda5A/sFB9cbbFbnXE8eEjmLwtumCi3GCHi5wtWvc0R1byJaZ9ZRczONb94JFpLj
8MxRA7PP8FtdxWJaPIpGwQh5uo7TnYEJtx5sM1T5pYdvmZfkj1Wy6+xYXwh9DhqFRByPcgqpuFgp
40JbJr2lIbghC53wh5E1e5wtiWgP8TxFGhQ9w9knMEUF+h7i+X56E5D/gJtNTPCX8ty/gE/R3UUc
V9amf0XLZvRQTL1NyZgOUFPsTK9PDVGQTqs6hvhdIZBDWxcQzXScQFss4rNuSbrmpn1ujdR/nwda
Vke0vUqsIJLOiOeZ8qYNY9RJBFkH03ssPJkud9sTQTgNKFN4rzzxy9svt+joiD/atfe518EUpH6+
j7lM5S4McLEjXdWE0pT3/MSar8ODQJr92b2oIAGiquOnrTvcGrKmmahCkCOIg/vWippcuL56tlM0
r1vrzRXKTdKmA5nzkWPUElQB3soMrT7jfP78YABbsl4HOwXmRZ7Jdc/nhGFd1fZh4WbeXjxBqeMg
ThoYd2oCpCvVJ0r0SPeFA6IQS4v81VtVDPuVo3QAhbEBXwrn/aZA1c1Y6EjpS7q4WQRmT4FIAJBg
UWadNyoKfun15ei6/0KXdrx+H+IpUY5iA1WKvHkeJi4c++XyxTt9cbhGXVP3rWP79laHgrHIO4UG
td4ZeIFJqro5o7VMhK71KxKbslNy1bJ/xtseRazuO6q+mIUKz/vuexL9b8hGf1RRTIkv6M+2LeYP
HFQBjUk7phqcFtiZWFTpSSVxuGHSUx4V6tpi1hwggH4FbT7TexoiLAuDAGpUYfYTc3eVsw4BI50S
5vDZdny1pmMvEfCqwo2zadHxuV3NUzJNEzQP4EYWNnd4SPfwJfKoCbkRLXWqbFde/5RLdSbuEuTY
Onn+YQMkPrSWfSwa4ELeaNQRjBz4L5Eoe+vnUuY9Fwj9Pq2FHx6flCPLGqVXOplcfrGdOVQWvf1n
McUSAa7/6RKE++HlLA3zEkWfDr/OEmg4gpJikMG1ao+lHUUrvT+PbpItuWQt15NaiRaVp0xcz6Vk
kSV7x0wQEpyhZzLO6lNbIUQDmPmRgNTJi46Wu8xfublkkJ/5/ZEEh1ZJ8UFuotbLERh7Xv1i2w9v
L64dTph6SQrmAa0yhbq0FIS5VrYmkbSH8sVg2lUnApod4taCnjKYnXQL+BwAJfnu7G68MsHd5kPw
ex9Pw/qEmP3Sv8LojenllY5Mov656AyhJqNPJ37A0C90IZa9NT4VoA2HfjuZd0+ICU3W1BAU7+JW
iPGeYQ0Z3eJJzESAwuL/YSnzXEsPkX1k2eu64X01gH3WPEW3m9qOVfUnfnLXQ7oDUPH5SiZiHycX
TVB/jXVaNkvJF4WNg4QS9A5BunIrisN52EwxJWzH54ImdkTAMhcAquBG92NWz9lEFMhB9Cp/1voC
0Jtc/IHJUe6Ie5Ml0TH/1vCs9SmhlGeJQHiCosXg9POlANBEidDY3ja5ndExHkSSio9sVvyoC74f
YCMqGGqToSGwKSKMruRciI5cMXBkV8jD0PZdp5odGv8cW9jI6q0pPSuulqQ9mW9zZvZ4XDo7nMjA
e1MVnDq/5jqqFVOz5ObRojfOtoFhDLY9AnJjifs116nOXaErcbhIuzWJlAAun0h1/T9wKWp67l4n
v1wasELOLH6qlkRLcsmCAh2rDnTcoSm9iq1e/3WCr/QFxZJuRqtx0rYCYig3dQpkzC+YgbDpGzum
qE6waUeBHre5jS3d12iMKSDI6fl4V6iP2+w2N3TQeQx6Io/aKNcMq17ZOz0AE3/EZYbuMCTkST9I
/foQ4SF3S0g+F2MRF1blQQQV8LLU5GlVL0H1eN/4REi+nZdEc0dUHr6NXqxIrAc0byogpkH+HmE5
e0vEMk+Qx759Rxcqn+gjnYsBQg7vnEIW9PoxAIjKBLn3FfO0QlKkoaBEAIruUHYfpoE8Wuj0pcaQ
6Z/3lkUPuC1fRbTbcU4unQNt2qsQVc8bF9lOjXhg2e7NDkTkU5SzEAaSDbMQPnbZxpvsECCuKa0Q
PwQRUF0k1vW8CTzQhGMFX7oXxsZoxGvycdBoKmMbTE99SoFIaGPSIdEI9bCcdikMIoJ2Onl9yFLI
GtRGBSgOVq064wbg/7ldS0cV5BqV3tQ2r+icZaA2U8QRcqSn5galpcuuFOVJQ4CPlOE7pDH309l7
J4CM283qhfKbh/WG+Hest7TmXXg1W3bvl+bAEM6WfbQfkJ5FL6s+IgPy6WMNRjiPQ5R9POyRQSyZ
hHwQgMK8t4CqcqKxh7MJ7uPK59KxIr/21C+wIAfpJJAjxtwShBIYLtSwKTzZY8cuPaEviwD5BSJp
1Jh6P14JqPCaewWdDcXRBb3OWGj7SyiYrOwMaZlMTlYu+e+8jRnPeeP9ijWtD90pW9ZDW4CsYlgt
3Q7MJfl0VShNBz+siMU5CxuVebp0cZt4TfPjK10JOIJDf0yEuLZgy0m0GpwiEhNLOvehP/6Gwq9d
DLLqcvdfj0p54YN1M50bCLtt+bLpBRpsj8tgKmJnj1LHKrPYdEXCffwgXL9OERZRljBctiEStRc7
yNAzRBm9BspD3s3OqYJI3oi0/ARkb2zsgyR7POHVY9tyS8KiMISPkS5kYwjlCP6dOBUtKTR9cBvD
h3IbqPTi4ScybNjwwgT/QcANiQxhPZF/ZsNfP6VortNYPWzlg7lu86Xma9+S1HO9APMDUZYrmYUo
5T+/AzNLW1pH7bBVimYNS8iWE1S4LV8T9dCBM6H2XZgjfFxwhBXdd5zjwfheBOZxpMrNJCZr/kpR
/HN0HupGeCJtUez/hg8V+FGLgdPpgTZwmh61miDSaOE3RoVVZa6VZ+cNyjofBXgD7d5fvIk7aLmv
vCKrS65PDNf6T3t2fzwHMPjFGGIP4dB6X41k5/jSjsFqCTiYS0Ld5APzBJIMl/PpZgve1OMhAz6y
9dRbUEtY0v2IoDSIxXKBxzX5nYM1sVnDJoSdoeZWNao9s0zVchz1q3B8PW+VHSqlylyHbY2rspjq
aEt89G5HBhB68vQbIBvmvoIqirpo7kn+8ylziNxBq4nifsWXieCOnjCg7zEdWON5ZqDjvftjxvs8
q6CR0nMMpOMVnlxJ1CrtBtl4zyXF86uAd/f5A0LNxoCu77eRAKkqWSup1wuOeyXTKiRz1vYMgXRM
e97xfe/V5kdTIi1bw4k6zR1ROuf5XRsMfkTBTtWpU2J30DaLhGE/yEhfXO2nnwVvrslIUNIScTSa
BNL68/KW0xE15YJYG+MPF37JvWgVnZgTQHL1L7cRcBcegiho7SfwyHxNcetyGBK32eZDdpXH2g/W
NJ8udaGZDM7jhdxV8NWa4wdvFVKthl0x3vRY9ERcukH/2Cd4rlzpH1NM+id8AiLBbjgtWLpEuvMV
lT+bRrU7nbQTpFa6Lsy2I6t7v+zQyRZD0l8mORwjzMWqZbTi0H5f7OH+zSwNhUvmTGJ6TCo/cVJa
PxuYpi9zzTcOx7wk9jqr8Dr5bljX1HrPaATIgFK3KXHhCnh3vpqSUujfsvIIBex+eUea6WmxXU6h
8ZFrOEkepvHfHE0vbMoSgX9+i+12+D4QAHOjg++MRVOOhlvzRoprUiCeAvCK7C6ro/iOz2n/dNtu
4Omjdmc782d3hGmlrWdJ1qOQU+SiGZiXVADdpAKMTXh87/1vaHw8XMYi82XAl+ZACgAul2kXBExX
72RNMP5YHXBS2m+wKMEY0r0W2+8jdJ/NER4riC9yLP3OkLI1RY2ZFFN2px7jWlfTQokK8HifZhKr
5GvGsL/g04/aNOowpXsFf9qh3M/icTkPQwTzBRj6Un8YW+v1TQtgUkSInzDyDtdprABIP0Nyx0k9
imorT9HTbrKyLTtatKM0E5TlpVjJ3CF7iQyj3wfGlNlpmQxYWuWgGZJX4kaCk98e9P1MwpePK69B
DOhJpL+q3xHqiu6DTIRsVBFSXZgaYRZuacRxQKufkRHeskY/ZxNC8t30RVVUAmZ/VOlXV8bHekSY
kq3nLOZcTzsWJaWy7H8HpOyPdufT19W+ziEgBkfzGHDzOCeRg8eSdzWr+d4uS4847F9+9xrTeZyw
/NOlZVSfxDR8mht2FhcjI6Qb6TqTedAWN4sRuQt4TE5YDhkqeaMegkYmYObZGzBBOtw4nL+9uZ1C
P1OK9oCD+iPOxIyuaT7vuc4JZn2/oncR5h69E3prmwq2yDUpQKWGeoF48hCaWsJUZPt15ahGdO/D
2HyIvtIFsfF94qZj8v34/429C5F1yzyZsp/qFKfLW1LJ1UiLeFpx+MMR+mFHpsF+STxau39I5xdY
wgT8uCqG8r4RbhyuWbuw1GrIUhZSjOYkq6uVMfw1zAUVAErjbc952OTC++Jmgp97BMtPuygyG6/H
ymzc+dj5hT94/6I+ZwI2wr1G4GQ8VjOBEAMvMyUphLtlvxTa2r9ZkHCNIVdZcUIhn7ynZIbZmCw8
8yeSOcyla6OwHnmT7Z+5M+Evd2bu2951qIhK75t3v2qvZZ8io6ebOiZYj/ICJz53lAGWyU5LW+Cq
TIJFXi/Oeh3KN4bx75hKGmtajVkC7EanruQ4UMS7PLmtc3yXbswQk2tQKh+lWJDChjA/Q4Zaq73B
y5tNiSZPjytchQF+3csuRc+3HHYUf6h3rBL0IvPWcjAQS3be0t9XZWeqvUOooqvTG+67bNzBmJ1C
zgTJwolYm7weOe83XeylXw7RKkYX7/6KeOTRjg8MPFFrPwPoVB6wM4/MGG3/fF7qFRAeqEfyeGjh
6PgZ08AY+AVAqUOMjytIPpUSfa4yAEdcIpqSQV987wTUMVWv6QJ0DsZG5E2UsIqbqRqzRLfd27h0
Uaqlg9EWX61wJXRHp7mBvp9b5S19790kY+XZUZ6o/2ZA4JbRj6DlyWscyjtxjg4Y/XhwNkixlum2
zT5buHZ0tCfWzB9u4QWWrEHpUkt4he1lYYhSYAwSldAqCxtFFniHkubxIoEpPGtvMZRDSKm2nS3b
FT7/UN5xe9lkb+yvLEjTcNNd9wtXsIU0v6NzhjtrQ/Jhh/45vmrjnXkP/AoZ1sTye2iP+rv0sT6r
WsyDl+krDaDExew/+m6KVi2yO3bdonl5xlOL7XjeA59zZzq1fyq+TkSdJb3PqwyEW0zrL7qzq04p
wpvXW3af7YCMdPy9bgr2RNp2yvopGDR4HvqYWonjjph4iwEVPE2PePPI8/vH+8SSFK3bgPmTlVw1
uPXdmGMjASEYKVeG/2zmyUMj5JC3rDT6TkLPaXijov1B3Sjw+6yFFuxoK0qGPK7MOPEIgUiQTE7q
CSaBoRY7ORsqgwdWQdRBy/I/6n7MsLeGzLXG2YIYbo4uDm2Ebsh20ZBIWrtqwZILvmKOD/W9ZItF
zU9Qu1nwysxkDFmBGXbfnVo3frSxVtUNzPfcOjut0fzGRCEt0xDrgus5NuEmF91G55LuJ4YgJoSr
ce/IqPqpSpaNKuHIwBSNYBhpFaDQ4YX01H0JK8s768Q7U5zPerznzLRnP7XM0sfmQiBgd7d8bOuh
dRevdWM8krz7r5VJZuKC7UjDElhAQ4D6AyTuZkyUstV3b7PC7y/QXTHMZMSknilKWbvXtQCNVc5d
s0S4lIhevV2Rgs+wryoSlUI38ETEiNkgbgiiPoxh7k+UfXurALO63MEwjD7izGVSdk/ZqliknO6Z
AhpnV1SpWn03SUn8mQdFyYM1kf7eU0y6oAq0t0kZ4w+1M/12yNI2NUlhFlN3Ikwg4W8daxvCJabf
ubGOFYgryeEYjbk05p6fUohIhg7djKOhA6NZBpMzL/aCfdiVR2VTfWX/pGa0fW74HkkHqf9WRf91
YUGux+8zbwhbptUBZ237EidazBX447nBRuHM5fLbNDleeKOARDGdtwuQ8zWLzVqGhKJ5RmyeIG9N
/O9yT8D904qfurM2xGSSBBszWMQec4iqqKF9HODvyjwJzN9CYdTQq1UkOEy6CYl5HpP2M8B3Zb+G
T540j/WbK6VQxW8oYAyAZyCgkS96Ra6iWBC0DWAzdvA+wEXj6bOieJUTP7q1OV14zPjLh1Dk3H4c
1H82hSko5bTFXlxnTdc1Mac3+GnBWand/Vpr9r+qIkkjPZMrDVv0rpXzO0lN/pQTgyKpPR840/R8
Pjnr4XR2mRDJXZdv71D7OVZf7LE6dqhw5dtdLiBLtSfeHJgz/FwZG9sSVu7IyjlmqVI/CZ5okO95
21zmY6l+YBP+DJU2C5B3uHIb3ZRWWnHujmAX4oMO41QVr+rhUtUbt4g/pjiu1Ntdt7MSIDVaokfD
+p16YeANG06okk4sYy1L2DyM3zESthITeXZpog2RebH5UhCEyDpU9mSk7NW8EhjEcpTKJVegrM+D
qCtzq3/n2rOsWA+WmlGK4yygl0LVYphWzM+OrjxSJ7CWAf+KH7xlBmlWMOGodmk3TGXMfjvdUP7r
8Q+GT9NLfMdKDFYTGb6pyledIHPJj3HFoJ7VszdLDjKohIp0kilLn+4BdzoHyWEe8RPWDZVqh4A3
8WRE4z6eMoHtFpZFv/ZqqgFpTGDGkqgzcjthGx8SX/bC54W2ikFnPeei4QzxBKhFrqXZeLpH983p
O4ydM/r8NTghRspH8pVdVyWYL6lA+/vtEAWKKkcHqD1dTQxWwF3McXeJrO+3VhS06mqDjEg6WkyY
JZDhnha8yOTdsqzJfjK3/B8rUexFfqqtqe80QxJxwrcNx+MZWDNtOT+FRFnxjnEeMkYRX5gC8T3Z
DU/gsNcQiBRaoow/8MbI33X/ULoE4k9TjjLJ/VTZXseuo65wWThkhRnUOch3T77dJLBeeTXLyfR8
SFBqIYp4928hsnOfUWByYNg+QI0DKpCXecfMwN7K+ips3hxGsshczDFADUDe+O37WKDbPME0k1Zf
BgDW+KFoSznRhgHymtbwGZxDCgBJ/kPSy3YPLpcL8sublkgoWvirI1/ylHzPn1ST3XTZ4ZoXTXt/
ftoqwDuv+zg025kLlExSZ5eFC0CpZ4A0dVkW2n6oEvs629nwf9FYhKWH44tXFDH8QklNTsh1cv/2
ajJAG2sly0Qfun7td7ViTN2vXBrsE3Jqxi98Y6m5Cb29+SFqsdXJMPVvqh2NlQmcYGAjPosYEhKI
h3W+DSSn/AnPlTUAfcXBQelFO1mbp70CswgzmjwybuMXO1+W2FWks12+jN20Kp70BOoOQj+/6eP1
AOBgp6jSWA9EHRxSalr+kS6TZpYRmLnjsTfjulZ9xFm6YDouOoB1acVi7qMioVfxlRLhe3g1Xzw0
EEOlebQ9cB/mMbiLjBEWZnL9F6gvSRuwXNyvqTso7twl9HmUBwzhLM+xT0IXRzclQQSWp7fDUHDX
0mA04+1Czv73PBQsA978ke9PRGCTxz0iFHpV8ze6JtwHoqygCoE6mW3A1jhLF9/e2o4vk04famqr
ZACqcKCwgTJf3OKudj7mVNkTh4WDRygbdXPXuDX9TDFyVC7vAB+XgCOOhTLt8EBpG0jf/XqbWBhN
tKzLr3DE9h3PgGAA3oRWRKdJ5Q8jGk6IxtVDlAEwGSnbBM/IsJ3gpGVLhMrB9WSGZXqbs6P0Mv5T
lMeIKpQpt1/wvQ+gOi46WYe7z/xg3J/1c5RDVowM/beWJVy/ZHhyl2hXeZ2V/MUbNefCOvgM1vv3
2xqbn7ZakxxbCNPfTGp59TvvA2vXpz41+/yOJbb8mjer6YKEkpp3E0V2DjwkFPsX0FhquN0dw3jb
WZrrMfMo67egc/xqHeHfpLt5+WbchmYdlQk91SNBknqV0mbgap9FVvTCd5O4xUKRkrDsE6ToHzSj
/Eg1cx1qCbCsdIneJYkSID7r8Wc+6qlG2rw4aYlTB0DQSTFtnZLtWVFf86MvvhfCcT88HwfkOp92
b3cqvi2REtO3HMFs3hWm7d84yGsFdBUISTD7wfM2JIvBG/h1l7geAZvKKUuUPr6ZrX8HP6ZzgDJI
Rv269G2kUq9NSSm0LdjeiaG4WnV/uBuhWMPNuKfqS0wkmHQjPiwfQ7d4CFmBzlenscgoBV5kzkvr
jfcUeSC91ay+NPG8IkNGP8SqVHjIZwXq0LZRnQO89bvScXw0mvwvbf60RWopfogshtoGu3hix6TR
MhghjaBb4cKLB8VXrZSsUwkHoTa+3buySrMtrAa+fe/woxcIaNxPPyimfScjN0wMvig0Wgw7qSro
6Lwu3hATULSGZQZAnwxruH5PIXc3jHA580CJt+3kose5cRM66O12qgO5vBwMgZAv7rlEuM+MFnrR
BzVVZq16/ujX+WaTEcKYCKMKxIAocA7F5raz7aZ0d52110BPzPe1oNTIT4aVy5UhOP/vLxE4zNru
7J5MnpdgMFOnQYwE3+0zFP8RzksGlLtJIC/b1N9mAAJ445yBEAhDxsI7VpZtdGfS1L1EsghVL1AS
LnOmBihaAuBE+g3nn7osDTMYiOYZkPpABs/6UE5j8KwoHr5so34WzKKkhHNYpCXwxvtL95+CliEk
XN8I48O+fKfiZ75dwlhVgHn5c95ZLwFP/4NbTSihNLOxJeIXOTzMiPO2EW5Tu3pft+/SYolmFx8m
Zofv4FFlZqgNAJOndJhPzGeAgTqWjyZomRgCatRl7aH3Wg2y2g/072b69M9ubQEM3/ihQQuHxFvn
4RRhkCPOL22H3CFsI96t2+Vs5wto+4sBPJf/HgjVjwhfwQpCKSOHEa/HgFMWlkMgvuKQjyG4tEol
7/zsr8cVf4y2ffy7dfQqAOJmxPybC/o8LLbkHDCiQBUso5ruEOx3xAUKDC0DDPu3LaCvaFCTPO7E
hnGy7pd9SLn2A/OeUxFLVWRpYUfCXjKxiYb03sdkDE/b0BPdXS//Lza4YG9VKJNAEkiMjhftMhkA
3rXL6O6FlxNrfOdOqALXzw3VIAzdbYVsH0D3Gat43IAbdL1SomfrCgh8ezb3BfN7ccFib5MfdywS
pZpb1OP3Bnz2hqoA4OFAn/sPlhhymDawuo11jZaFDQY4n6x6JWZAPqNOo7bshFGKb/JCiZPiJe/B
savvkyRkDaFQc8jK0mA9y3oWnSfDgEy/NO2LV9nvFKZoLH/awV9tOWlVr3mVuZnxj0qdvXn5sWWW
1+fJA6zv1TkWywAucxaDTmwWFL+M1zcgu6cvb9nBbBNHIqrDZzoz62Ge5xSPWk6jz4V1F4MZ3HIe
sanU070GDQ3/Rhf+gcmx6CB9DcgNa8JsIKN0OS8aaydilDONEJTj8PQ1fRL2dHG4jErjgBdmbqjq
sYoqQ6ogyzXGjVmqNVehUXiqZZv8827l1LovWr+qIBtz1gU0SWEsFudpJFQvRuIPqzV+9O7gFaAD
ctRUJDG82L15b0xaCPBfw+E7ymXqog0PqaRhS/LNOBGSDEtPrArgd8o1pRW+1l+8yrZK58yIKUNb
x+eZjpriWPf8QnUj+rtBYRiditiEjSzB/pPOYytBfoAeO4kZK/Znhx7elzJUKh5QVNZCyllL7daK
a0QT6SQnu5KA2nuGrIz2AtT5wlWtJgRKGBC4TVIBobPSApHBsDFAAdnULSJ274uyDtdhTtUbkw75
RDuRcYyTtCYVfjbvNp2T73lIEa+V/2aoX2n0Imjszdb4EVcx3XJnzmpMrtqpFdrIMAhxqMxO+/08
LjytKGC7B5DLALpJ9WkMFm/hfeTWJc9PfSLssxOlNykq4g6WKAyY2sU6989RvnpOH6GYOU4d0pI1
8j4Lr77HosmyVnIPfMA/JLaEO24ao4+3S/WcAYYJLN7Wr34ABab3TO4cgiEg1U8/UhTt+D/oLefv
fOwwqjntRheLULV6wVlesV2KDP/g5PvVtQaAX3U4GSykqm0AbZaflEV3w5ACd6gK2s6FsNEd5L+5
ulfNSXojVE/xEq5immjmxZrLnbpBgO47udTqOdDjTzRwC90EX+KJJ9araKd+lt4SJitfELO1i6fW
TUY3C4AGwjxBHgv+0DyjtoIEsLfK9u7KsHo5m2Y7sry5uYgHvMxFOxHCc6zbPkB6qXon6yFsso7h
wJ3+dDJQ/zmxoKyZhFSr1UcC1aH38kXkgqX2J4z+H9Jd9z4CODMoiHWQFNy8xMmGRa7F9VbMgMhH
upIyN8ykSkuYOdc09JTCDUnUKZCUnuMd6RyJB0gzwub2Pr+pt6gIqn9VBrxq+eUd7HtVyHRtuzqJ
iX90/s6A1uLBzpWIGnBhP+VGsel5i2GIsOy+kPfFT1mx6XSl/CJL1ZbOpHtXh4n1KTINuQd76Yz2
lfGP+HAh8oWcwUcp/bsHc71JcU746YyPmNQdoSJPtPDX4kN/xjoAXzSs4AWSPhboE7b7E1B9vrHE
ejO6lLHHGLnEZY8pIPQguSaRUwu2dPm4zFJJylvd4TxYBfSzRtOGLCHjCDAdkqQt/IJOPBXTazyM
vaX8sF6+xpntv5obGgeVzVXeLOSfh8BVPkLj+jvu11S+1/AYfyFmb4baDdQ4SDUBdPnJ7NQ6CnkR
52/Ob8a1UzYx6usGogSTw+NymS22HcE+D4+fqLBUz08Y7yTvBgIbaLB5typMgq8iO+Yz3p6g4R77
795TbXyWRzK4y8X83+GwJZBQ8GqnsdcVIXymQRPFBkzhYWsxj0QiLirnt5Pu1a4EIOHYqJMVEgTo
P+4zbBa2BPtHo3Q+8auX4hbYeB+d8EYYj5tT1BJQiccyU3mrsjruIZ6psUK6IWTRLFEyMtWwehGb
0NjjMzshemi05TOqJ+SPSb26+kosPIWTbAQl0Ir2xrJqudPYHpdJczT53NggkSqB59/aBuQTyL+t
+bHEJVZ3W3KtF5wqbrRN5azWhJYX8wva877zW/k4Fg6T8+dLrTMZCgMFuUxNl7YwxFM2g++pSAgi
d2g4WVwg8Eis0nYyGtRUTGgOZ5OgA6kY4Wg4L6/zA40bOdMYVgYk0qap8ZxIZi72z67BgbTckhEO
J4vw5VUhELUCpNFRNLjYI/+8tyXH0TYL0kxIlwOTWQqZhQFfIhuZDHJFrr7JeeosvGP9kGeOqNg6
s7GnoN+l8WWoFVg0wukprzkhoAFdSItjeGMPvUXuGpgsLFdMhChMkj12VVhP+nzk51mcgI7EvY/a
re678pZhvZw0sDWbpahLQfFq/nelqd4XbQOOdiuaGhWogM0mR2auJfmGjh0UgyKeJgZ4I5g4kfz6
bogGWh3NLQDaCp0XMkDWimza20TlNJQMa3iRgxcVfYR5uKM5IikqnTTCDczuBiyJLQHQgF2piKgF
131AeJwdIYuom3r5Y3lk1vjI5nh0W0zNrpiH5v/v05dlshBMjPHcOVQgGkOMBTIy/MlJWJs1wRTQ
0AgW5fjGzwN3bBKKy7lIfUoPmbgnf4K8ACA+tosndlXaSHPQb3FCXAr8/Na/777bt3Zdz8pMyz8b
X+tR+dIQ0cUFY+jfK3TFG+rX3RNmG+cNijGsk/N1/rhe1rx7/bDVzbUgO/Ws8x+q6sI2XDzT4wz3
fkrYuYup8MYUZITWUoWJ542xTIhDp1ziYHQPl100FaUqXg6FbJSrzjqeOaBT1JBOVhvBG6TyAgFh
t6K2iOoEEoU8UqcWFm/JRyPu/MOvvYpubyQdC73dckjIDpJZMz6OK0Lu6mQQu0HrbJiX+bYO5bDz
rw2HLqNecdnZWwyRWAoxY1+7o1jpf2J5LxDvZweYTG8ZZ0cnlhdSHmcfnD//Q13RAT/+7wsaIQ+i
KSNJy2OFXR+ck5ah1R9sDsakCxtpF1AH/UpzS4bSJ2CKX52w9YKddgwYVuHNEIKiDDH3UTmOcWBf
HkvM9vVH1y3w2EkQMLusDml4wZf/qZ/9U+XJoL5GXnOBujqAXP/AFqbNwh0qGBEH3kl7BNe4hf9A
d4NKjX2CHJP+hph+4ylQqAPrYSW3tGpNMqQZy+OAvI1Huys1qSfwDOXVQkxSrvrQJjj59MUCcHic
qNya2IODlYiz6aMlQKwv5jvwNZY2kUZvo18WtFhmYLsQ9L/5oPLP5QlCrqKYhTXBWpfnGA6q5uVW
MfUs8F2NZSLEnB56KrCzVdLXBb11dU1CSuWe68nbqYPuIUUhWDjRsyMXDC7ozreAxXAtvfvpC+wr
2bXazBPoMn0OhvwwznNn62I6TToazo7MdcqN9mQxEK5FBhYW+XCQ3A29WZiSjNrhcM3aEMORi4Fq
fOvyXVG2U9pmgcKUsVs0jz1I8thNjkW7WG3UWSbFKSLiJhmRdDc4oUfJ43StrFYhKsZx+kvCE1ib
lo0o9dAXG3lTSSepznOG/WKwiXDZjXXuhEwNTWWZxeCgPC5AeDE9qzH3StW5WgJc6laGnmbhRUAs
MuNTjxBFbA218KJCdAJXYCuilIm9m4wMN3gFauxiGAbvFC1MZO4yNdVIFWw4Ir6uI5rKOKyARq4R
7GrqaSbVwEhuFBshAKVC43D1uN3/HAAAbGKB7RXI0/4kPHtnuYkaom2nKvW7Zs65YSpSrwAeFT6O
5EqxE3DHzHCHd6IAbkw8XxIZyMV/HBa+ARIymmb1M/e3xWMi1/NfJ9y3boxgXOMKU2VbQt2fXaWP
8wKQiZkeLodtfWOSUsU5rv82KbHf2DPiPzf8wkUXf7fw/qleVdVVOAjnC/X37eF5D/I1N3aC0C2R
fuAOE6wy8zbmDPF6K8Z4V061oexdI33tHMwizBkBrGHL4L6RDsDX5fcsEoH7FLCJ5rmQbj8Ckzmz
mHGWsLjC9c8UCSZQ/qsYFo4cyquhvJN11y0IknUoMOVxATBbuvyraWLNtWQwwAIla54NFwc3YM87
1/jRVn8WfWceAXO6pgEWKM07VdI0X1vBDMAUtw4fyfaB4IPnB/R4F4e1o809eEf9OCygC3P7tezP
wF/8Vso4oz5nqS3Fmbkbe9tbUzPHVoAgGxu3/3j1qntzVH2vlUR4N4MttgxuvZHVe1+VGgST8INx
L4OjdAd+iFyLT7rMGBA5S7KIJKRRdJD6Ryz9ULCqEcKhRU5QEcp+RH4BlNEnVD3kV4/r1cK+u6xU
U5zqa7PyPXPqFK2HdA+3TXgYTMlm9JeQ48zvKlSbd2NS3QpU22tRDSuvYxM5bxinPjC7uhwUY11z
Su+70Ptyu0oizQ1ltLTSr2gLWrCDIu+5EV2UKYLjpGk8ygOXLL705VNrwCIx37Wx2JX1hfCRksA7
1ZBVmx6SIUsEvPm8Il6AXG6RWuyPqRqWGIL26w6/r6ltqRB/DHTVTGwdyLO5w8PJf7OoSgBRS8pe
Du7fxAjIpMzYgbKxTpAJ+5UWSsxtJ4RRXLaEehMuOT1q4yoR7uB22lvHkBl5jUOdeyuvkZdpRqhG
DWUQLeXmkqmtIZDn/S5pySY0gUsG4LVEGyY0TBUA3xWFwyxo0CA23sAxw7blDfAW/MR2h5vNiO2p
wLCFkQAk7EMKpzkVvyeHTGUBDFnTfwPNj9+ZJhBiYClaDat3mOJjDa/nrG9j3Jltr8lPbBk5wBqy
x8fDr7gDyD1NoHgYQBKp4B3tAv2OaGOtoY+5XaCg83+n5jIAZFzx+NAWUZklgdFG37Ohx0OjoyEU
xk3m3O1Vki2sOePjb34cOPscDxLpc8dPYwlPkIJqxMs2obC9hJ2YLDViXW8opleWz855Ke9eWQxF
tIvNneNwxUax22Vcxts/cqI/uHN6NeCifXOYBi3cHqvzEVxHfqvsKxXTO08LfssOd1q0B21ZwU7Y
v5ilGH9FU0oyH6FO0SnXiuCh0QoC3TfIM2MgYz7knE3NVpIoeh/zEQNU5Wuge5k5wsTCahK3+3rg
suNedQwvXm6Q3KJRSC5n7U9BsP0PrRAzv7seyavQaIZb2+URVkN/lyISKKXzMzAG/czK4V/HCXBE
GWP7e7WULCFVBh/0rXrQ3KXc9jCC6ZEDcVQeC4Nxgn4Yn7Q9rzsSBn9Cw6xSB+dKN8DoF2vFd6E/
fgKCl8qBLWd9dasH4r12MwxSIxC1D/+QwaMWDS/dKTbJvh9WUGNcDaqs1xGwoKqjpcVV6wKoxBI7
P9SSSXjvQI7GwQ2GnYtcB4/fN84yiE7KUpdIRRDLMj4s9YZ/7DfQPzSBudPFL/joLPAyZLhyEWyJ
1TvUMggIKHe5fZPfER7UTpwIXaqdgYv4ji41IQkWZ+JD2ysQn3j+CRmHinnTDpbqr0RiXRyLa8Ki
/u3cHwEEfurJ18/I+HNB8rscQIzlNn9CuMiQWVryfB/Q7dvk4VO+cp7DVEE5rZnDqZx18/wBUMWI
yj5UMiPjfFuFYDKxVHdLScpdwxqqBZ2+/lI7C+Av4BAlOhtlqMy6+JBvoBFtlZ+IoOfhEJuMhDg/
yJaDTMTsdGunnhbWE4MyWWsw9/PuuK7czNaScWbx/MFsTXxmdz+P8n60pi/OZd+dbALvwW+Jd0nh
oF50uKylh8uUMfkI36LobvXhHTGjUY7Sr9DNPBS2gtapgKBiQU/EnDhU+rojM5Pet/nziaLCFMLy
0sMsZmdM6QmaXcmB3hJp8qlEoN1NqZLaCFXfqHDjoEykdgme/NSneegCeyD+bNpAurN8gS7ZLfd6
zRiHRoCru3jOX6dj8yupcnWcjnsYA0hKTXdBedsAVjhjKTxrrmprgpAeEDLNSOXgSDnmnBzJJySZ
onXgbJe63D5Az+nxc5YvL/oextxwqrbobasov9tk58/GgroUgwLOfEqKTu+m1h0qBHpy7o5wQGNd
CXEhWbB5k0SZ4w3LeRplk0/wWMYdB9PolAUmcymYmT/RBYGelQ1wQj4eWQIkR0KHyfaU6CLFddzH
Syju5oM74hYspTOeKA/5sGAkfdUq5DB/p0fJK8MoKQ+L6GHmBF6AzaIL0INyHCy96vNZKwNXwHVK
/wx3jdPfGDGt4iOxnCfDotdTLaoybvXF8I6hE6nQKQqzswq6/oO8xwwAoud9b3vj88UbS7+qoY6u
z78e70p1rOw/ctijTr9vAbexOxhsoqqdjigrJxO0sPfkEzn9dLXFzRwg3c1PcSEupja6MXDo2QX6
JtiGxkRNdkbIxrJS7XjHXf+Q2HcwxPta4JyO+agEcRfcyflLEGHHT5aRquhxcBnTQrT4n89ne1Z4
int5AAWvwSrcV/xC7Umqbj94bI0S9j0JelYm7nXhYTlUPtmz1CecsnvOx1d8yUVo4H5e3wo/Wfc6
39rKD1q+oBjCpdvS0nuGQ9vUMJUzuq6xlx1HI9kU2POZ62Q5HLe2qYCHsQCxh1Fjd7VSQzGPn/Az
VWifIzcaNucBU8SfYJz+Na2Wxw5rQRPABYsAFiEa9NjPWeLmgzpxNLrpnj6M4jjFdClVtd14iaQt
sSh9SuA3MsoiM5s3EHrQjcZl4BSe2PiXn00eYPq/Qxyrh5qr1XKawOaKfyL2GXmzXwDk8+46XwiJ
LMWTlCBYo56gHCIsb7Qbo6v4/aC0z6XXBbhuHQmyVmR0LObD5YwHK/ttSZapzgwM4nQ1g/f7WxTD
eqbcc5eExdlKVvbCoQ6FnzLaflTKKJQUkY6FBOpWwI9HC6uPo/Ic+87sjNcuvJcszYXiMSXyljUZ
SaEWyQQ3tEwEymNfch1Yyv5qsNsw08XnNrQ6/KHHpSbxO4qE3AwH5xZuT7BoIVBcNJL7OFalSaEm
UP/8U1xeEf/Y9gu4QS8fQSLubgMh5ftYgTdTejurEju8WQawPtuiR2Ku8DW6DtPVJ+6mT5AicC1O
m77Ga/emfTJ6SA7UIzlXN9ao/d9AFWKrGcjHP9xTNeeT+meWMvt7pYV71BXGdj4OF6TRXkFvRI58
rdZ22boDZC6nxDjSRMmgwc+415us4uvbqnArImHpaponvY7GhhoCgxm46DD3OTN+/s5G5ZGVySJo
0NEMb108i5JRwuk6xWe9GCCoWjSC4NfzBS1xFJopPCJPsc54lZjcWW1T+12ABjtbPAnCkHxJq0q+
l7/W5wk98tQQkL5mhd/NGn6fgAwczCy3AAZ/ThwnNqM9JEwoa+y6UzISlxo2Ioi6LFDIKJSdKKpR
izsl8Hr6GVtHJ9LS5yonx8l/X5HbAng2FKNnziWubWpx03OQI1Bp58YARgJ4v5lfm3ZySiyLSAe2
+MkGFqyaJj4qzNCLTwkeZTpZ8NqBRpa9eRy9WhaXqCRnh2mnC/vnnw+ChN/kZdvWYagm1DkzA4gQ
y1R4nJ/urz7bb0k3iOAoA5IvnWo3J/PiaBvU21N2w/0betoiztYmC80HVtokU+wdrPvhwqKlz73q
BZ4SBxHELbF35o8PZ4fNtyaNhfUPoyCiqRQJ0Md4AQFbmctqYjPNhp/rUTnxjNHROe6lffrLeP2D
d/8pWDo5YFpRqKH5+PlGDhSq6tU9QLf26/U0CVDE48osHpbgqYTnllelhSWVLayNOBncOdRe9dOr
93kkEQOlVk7hn4fp8DOeAasgCVzF7BK1aK1arIvkkuECN++NB3KRg8We1saaeN7H3SgEv5VnZvUB
mTbPMlGcQGIX+1EUgPSL06B0WoQIEqhcX7CWcDilPhFmKHiQR/S1JsA/JGZJkTzUXAiigaDsXuHg
rmxezishJwkC1W7q1Lxk4eyCdgqh8cBOGaewvsaR92YY9qgYFqS6EaCq9cNAb9LAsTSZDTQQPfG0
iTyzXEaa3fxVDaokfaQ+YC+zS4OyNAHglIhQ38CODL2pKtMLbGdMQkPR6Pgb56f4UMezz6v1sm5J
G55FWcDxFtakm1heuXEtETCG2xVunJXjOxzkQXuPrsXfz0wHM9jvIRgD6G4Wztdk9JtGEq28/gsX
PJ1DoYYII61rTK8DbYkOPAYDeTqVXvo2XKDLlqPd9KLwlYa5F3wmf5A0Juws2UkRHr/+HytUF3Im
slRr9NZazddRVoMEDHf8ZHdXIE8ov7QKjajDHI+Z2Bm8n/jts64i647NVqXXfGSOYQJa8j8BvPPo
dcwr3mNE20RGeq2IinulxrHDmqY0ndMmtRq0Yg34DmN835NTN96U6Jdvk3T++OeMv7soYikqZ5qc
U8xwCAeHIjNbxFGG3Q2O7/KGhHArbZprT3J9NLKW9TmjltBOtnU8RUPLgRznIq0hmzsBWKieHv5C
YNiFajXHkpgnqbSJF8qgAMYXqPMNw5oLvIdlme9gYiILUEbvvl9dk4MOeKYWVm+jqm94IGts6pFh
4VvDVIyZDMOR3kPpRpB3pLAiCwJPELpdUemOpQmFj8raFWT5M3eNqglKeqBp7IjmuQgPNjk6N2PT
+fbYqR8hLWPl29jJInGIq0TmUP4Cf+vasV74fXO9zHtiYHwdxv1IdU/WZEtQcxyR05sDw8Dlz+w0
Y6plxFOWnveaxa2SOyvkLJ+9NFOqd00YsVDBRngias6zRWTms8SyH8R2gneAtdwqC3hZDyH3A7gy
4N+BPV9DQj1JP4ZflqFr4BWF1z8i7JrCrbqIUcLpGnkjmQeSut0Ca+8Ve9E9Ezk4gh4Rrfo1JEvQ
9htzgD7ioWSrlkRwmLva8+Pg66D34a1W6aW6Jyk6+o1KuTtt3U9CIW/qaPgUBULXcgZYGqo28+hB
kcWAIN+dPIHz85J7reefLnSaYs0AbXnSEw1ncP5lNJdY+eDif5yd0aN2adVnkO/7Qhu+wf6TDDpo
f8EtD0bQo0PUZb2AL5bBRPyTqbIPbKzLkJvH5Rp4Sxqb2d5cKJNqIB8qMua7BkZJZrwouYfpEdOP
C/gI5N1MEFcGD6PtIj+HVY3Z7vCgvF0XmFWeyBL6E24xRQ+7awACir9ZrdlVqh4KyY253Ns+QqCD
+qGw5OiIDBKdngILV+5d0MlMuTy16iCFt+TdpQKMOt3E/iMUtm3auPqw6DKHOaZWdFs/T+2kxHXn
kUCoXzeymga0HzgZBLL/IJ7GicMBuXsmMaWx6z8UVW/ENOYX2yd8m+gqHtIjYULCdjRpFVN4OGM7
DEgWCnxIfO4rzQ+1F1zQaZ9kCCKppC3ff/mUEtbD/zAbF8SN1CBspNIK1mqOjTJsKVHg94KRAfKs
lGKSy+/ieGjM7ibyeY+rFZ4X5MSZiuXVhKV9c6jwx+3Bm1pC9Rne6Cf0c8XeI/x/bZUqRgYPo6X+
zPHoUV7mktqutpG6eivH6MmOnEnoSWtMUD7yaf5OQ2MepjAnPMI+73JXIg4zaIUClNZLXSDgfGiS
hymamIiUnTlwYrpX43vl+Pw1asbcHMyH5JmViBHjjjAI326DIO/D44GL/xUZwsy/6HCIMSS7D0/R
XCWgYif5Ul7Ubw7rDh2blJmksxzeeCvKYo/37rCS5hMPRNXyedcHUQ0yklWyh7fLWqJbdPJtzl0E
pJTHc0lSc7mtduJtCaPJA4Ei9DMTa/X2FZzuBxevXGen8KBrGvk2zDEisGr4dIUHFHa5MsMejOzq
edXdWXDN7dD14z6e8AnI+Sh2tK/x8jEsYytQGhOh6tzDLSzBn3lWYUEemPjkMFPcRPv+pXP8NFUf
O0vEFafGNgHPwP/HcJkS4TLyv11feuMIPB2/sRXRk+2sTPk6/U0zW7nAnoLaDFN4GZrixvWKZD8V
IsTyJg2CFU8envrrvtV2s4Q5ELZ/J5WPY/0A8kVYkXtqSGoLtTRvUuRVShVAPo6/p9YX47BoiFBH
Jz23q1iYPOkmpMfRdSYlRFIhecua1ootOzEcxYIrYtEE77zkdDxjKK0/Csl5UflIAFRKHsZ9n041
SYe1Jmohb2H2eUyM4+GgopvcWgvt1ug8fHsQTlQ9A9HhDSiK8u69G7Yj4NesJ/EKkrEx7n3G4/51
YD3PPd+eQnc7Njk4ticaPr4r8sV6eorQMs8CZqCtU0jdUTGm+ndO2c76gpo0OQDvEgawfvwCiaJw
STnkg3q/UQMXKiSEwg69hWbIakHZmn5GKmkbWPxB6dra19epPyDHbxEqmVyXQ7BbSz632YsF6Tiw
IIL6FIFi47L0IrEw0AtY8w93JjhvLrQQkkK+zD56TOnaaUSwfPFRYKnL2cGDPDA1IJaWUPAOzi33
fqQdGNxTKx9r3iv1Wl7FRqvarNM7tEY1b/cyymnaHp1M3sNz3tQVW661enCg8jkmScvf4EH45Jyz
hB92xofdZG674UDBgxOZwYutpuVnLK5K/mmILnnJoOsbOtZnASU8DcfxUN1mvA0ZwVPUHxAajhqN
6SzzbSr7kkPdA86tWAv0SEDxAOH3HC8apApD+Xk50sFK3IrwRLMcSv33Qv70SNJnnSlEDPChfMvs
8og2fpJWdcmylU7znLyLGh1vUwAe7XGSRttR6t29N43P9+WePVqcy4JynYPG6Dgl1lO7QDX4qk6A
15ARLF4usZ99RdW/nVVoiBmTsrHPxFnDsb7ixFkQa8X7xBMzxKAHtlhi0fb1x/16dRYbG3i1oXor
rho09Jh+mNvYJjWw7KI/J1A9w3Y3SX2xj7HStOfIxI3ejFae3sJqpl4nNOZ3RV8j9DwL1knW9dh5
1itcruXH+xJ0T94nWBeFkai9KGSK2AyHmqFj1vy6Tq/Q6Gtfu60I7uSbmvMVYY1THVcdhyrhmcb5
rLITPsBru/c9lDlJAMjxsbvPHvapKoaJIR01QAhxQAdRty5oIlYJjSdhCtoiK4QMAkNlLNiTOvNR
yf7MRK1eH0Q0aZSRbHZK8EZ1lrYCOGIdSzUjH2HoTgOty4c9i+HqWffintvfeyW2yP/YBTn0KTsF
6yp1S5LmolxrH6bqsIGmORwhhcCANjxtEqQ9CrgprPaxjI2uEjmwN45uXGnlVrarZ6eiVNArz+ij
qUBau7yiFo4rT7yN84qexzpoDLdNrvP+RmBkQLKKgjrCGFzlZ7gPOxt+9GO36N1JfDJx2uh2vW61
5+AD2rkEg4YjxWOBO8vENLmLMOh9MVzWbnyZyVB38jjO7FlpNP0QQnjEPLJ7yNH+xCgjWGNnrH5k
NrxsZJ6ANRjzBYrf93q5CU9zQv2i5QMHjKHfGyqFLIktW4e848EoMecurrS/o/1PTql2q47+h6t1
vlZwUTG69Wx+XSDq0kwOdh9XUlkyWUjuBIcrBA8TrjNQCQz4elLuxkH4QGQHnOwAel/yq1bhqxUo
IIEbbmw+jB4F/RqaCX7/a4CcDMv1u2zkJr9zHYa7mPoGZtVr1YbZ4IIfJI216N5XucK+ZVmRZCgy
y4FJ2xAZmvuzv6r+TEAn8OYqcNWjuTQSlGriW/+esKodmTW5VfJw/BMtdhJxUP+4VXBKdC9U0zU1
Y+RR+cN1kb2YQAf8chtQMk/2c9lWi4XRAjFUOCIfuOgE4La1/XGrAtE5mePXIDwG3bNujZ0CjJ5a
mq7wWuFRFZ4f24NQalUhNuSkLy2CdgcHeJaI7bIwUWaM8pr+fTyeavVmibxz0uBZf9922cAXMWJg
v719leHJP7J8WXhIwTexOEJ1wa5x7+RrbxdjWk+NLE+Sds3Quw+4rUKYpZMf48EpI5Jbm5AKLhog
PmRr+LNrreLeDEoworlZ/G39w2ChF3NLKFM48QHO3jv7B8RGdmzjNT0zj4X7QSXMNF+shKLRZkfH
y8/shacrWEjtuU1Yad5Hn/qJusCmkerKidf71ouHya7RHXaMeadawuEqSg0zLISNIR+iq+cCxItd
nTbCSx9QuOeFvDnli5+qHf6EyBThCtY68GQA+Qu6VrBtFUcvJCQH8obcjB+Lim7/1KMDRqv0GvX/
sO4sYnTPPZrjqQ4G7KZVrmSa0Hnn3vW9yQDHvSGglDo3Rs8uXjlYtXfbfLljFlXqK++C9qE1F4qp
fpawi4t7pt2EM6jm7BEpCIuPON0bbCmWVSN3KW2WfUKlhMDYajaaJx2jsEBbjPKlEL4UgGgo32Nn
D+kjwVA+viMlizzL7MlLooaN20UUvxPNmksOkE0YmwLVhqEwYhdanMc2kyY/1GXy/vDmTOY1H/Jd
EROc1G+bk/jAKCh90KB3Wt8k1w+CWV20ofRQr6Sygflg34i1T95zQ/MXVHMVVAs6DZ/RaRQufH0S
B/dG/SZbZDk2V9iZaRLPffUfhsx1/gzcfvEUTb4ADGZqCHUO7WhxpIylgVc4XY65SBzsdKjuH3cp
wyOiwV+lTsBnM+XJ988rki6mRjN/X1HIhpZLP/1tXVTW17C+Z797ezcQIUx0WW//gSuSsm5dfSvP
NGyuczthvkckU5B8TyLF7M4GH7yzZRMLq+eBZMw8uLX50+4ZnOeuYAKskqEgKt5UzDpJDPUjXNJE
fGVcRs05Tsh9LlCwz/ya8rSi0iJdPW5wcUU6rhIZT2l88jVCC0sPtRQJeoIPnl1r7Nt23Cux+AQe
4Q2VtHfcL41z/VgNdimZc6X4BqFGCAykyZ405P5CWGy1weSGDw4mnjeKFXYpq6yzQb8/GZ9LkbLa
8e96XCg451MMsIDJFeA0dWswxcznKE1jzLzf+5dBZhCSxOjnaZ9/x5GKqpmU1gR64Prmjzgjc4i/
z6bCJ/jPmiBjT/JAU4MlwnGJA2fIWbafQ8hAObiG2tXV2caA4h1v6eQOaJAacci6ZOpSxpzZWswg
yK1hV32jnUxZ12dc9LVQqgMlyvoNrBQbU8RUwjp5Jt/uSFWy2cvSK1hET9yTfstB9jT/RH1nGnVc
XFDYDwdC070erOkao1hxuNX3Du5z5M5hD+sSZhvFwdJGG1kEcRAt7g1Ii6tlx6NhiaHqHeNPUHX3
QGEQc8g5Uthe0cCTL/0YCqM3xEZ+V+F+nIGiJMSoAorwlqPcyN12DkJoM/zoI18lv3QI0Uw9JcAc
/QW3g+K0e66ssnM6z8ZNLhacJOp5te5OpEd/cLljb9wP6b5JFHAwbTgNLxfcHQCGasp6AnlByBRB
kINBTjDOTHHuBddw9Dx2SV490RYUSopfuA56z9S/QUZNX3RbmTeH6SeOXijiTkO58Ycfw/XRpp5T
EpES3QlZjbWVasCqwN66OPAqNsqD80DToh4tggNGQe+FI9I7OajqHCOWgBJ26X4YQYNiY6ZNXxS3
JqsKZ0zwKseLEu6qOcOAFA+jhKdOeK7aVx0XDtcoqwmOwnKTLgzNZWT95HlmNoRNZPeW5cD5qBSD
qD/9IKQ4Q0oGRCFnlxiJsHwOtRTilVB6rFOlih/jx9vRozqAe2g1g8t++guU2bDRla2bi9tKSZCz
Q1/68JjdX3wzsBXiXQCBPl1LYm6pMCoJ/BH3r+xNwxIyKSL58uwjBk8Ck4buhytP/yS0Ygexgstf
NQvJwGdRlHQ4NKD9aoUVkkpg9jOx8UCDm9Hj3pcOET+vrhi/hu/N0kH2JbYDbkvz0O3LdVhti2k3
aqHOyxdZF532sVe4K7B2iaIiF7VP8ftGfn8iWjHWBflcxETzJAyQ03MrPo/jKE/f3Pvs4XxkuWO2
5qKvdzp9m+PdXRQw5Px2Sq1GEGSC6r++KC42WcNHy/IQzPz3NqXQT1d1Sln3j1q5qbJNQFHurTn2
Hlml7NTFWd1adKb78pM87ptV57owQHbiIyBkRXprfMHgY9ZXfs90aiFcAND/2cTL8Kbh4iZhPjC0
uqPDfP3Vg5UuQzUKyUbAP6CxpjdV0QmLI4AWJv6dpyRtOKBR/s3p06s7ziJjkM5DRN/IZMCLAxh2
g4Ix8Q8wL+hIR5i35iTU6WcfjJOaXFBI7/l8lO+Ik2VqMMdHmLbtNJuxRut7U8UysbdsnoXKWEB0
6W2rcEybiK9qRo3LF4ako0x/IoL5S5cmxub7K9CAfldo0xjnkntZE7B8/FBBGIAp0qqeDjiD/tbO
d4ckD+zYKV64ROGJCRrPxryxZRAsZU3r+6cvDhw/sWnPKLBJPJcqTkt95SUUuOYAy5Pnq2sdBO4B
4gyACYD318Qjtj5UZRkNYkPN1B5MO//sfFCzyA0CCgtgUi3pEGjkvAkOnaa3c21ndJjbpt76rKX5
AwPGjASiQhrQXi9LLTBRjb/VFj30nKghdg6UWuAd8vwwOa5BsP7t1/detxpT5AYWjJZxm4UHO9sG
v8YiTJ1Ew/QGNYAjXRDWaTa0LdUK/H4oXXMjhRnxxNsVs8HJ/lBT4/GcXWgfhixgf/ckIORxVBRv
XHOmq5Q4/T1kfIIAjpoY6cajjge6LtNWM2xlY8TmMHkWN8EnA9ltJAL4W5RWmFaN9GGH67qgsknB
rDqWW7WLiAT7NWvEssbKnQbSFTitZdnp/1tbgEbDgks9cU1u7OGeQMndtJFZ9Mp55MThyiqT9TX5
0I5owkR4/m/wPJUUJTsIGiNbzHRlcfRGEZbtQEgeT3SZ4Nv+q1sshTsk0scWDVuHMn6xh8+qpbDW
gg9ZgTJ/XEMgB0qcnYcPsMH6ypUogV9MPCctImVb2Ygblboe8rilV49/BYYpscsjUbJcuk5pqumt
3MnNuq/chUeoMEAnln1XdvF6/bOlq/w4aF7NrmaZLR4Yij/nMxNCEoagvTdradbUQUgm8ii+Q6+J
cn/0nmXAjBUco7P3nbuJcC11A4/GEnrDJ7IiWY6qvBOpkpR/6YA1uqhjknQvZje3DkPq0QAvFqwL
keaDVYKqeA15cwYbEPsYodkvcutS5HcJq8woCjVWPo9MipQX22ez032MSHrW+Yem6OXCgQEQiJ1M
r0qKNcTuUsOB083Vvd0BLgo7sV4iLS+LqLpQI539zxHWnXVOio+My8O3CsBQLMEwj64u2rlCvu51
MMvbBfGWsaiK6Fzt9IUhQF3UHQ6Y3tgmhmDTcRdeUHjnsiqtXpQdnIQas/3H3LKRZ4UgtHy6p1dS
fylnnMYWaGhxbVXZUzxQkUf9G2FTZ+JBvfMkUTe8zNK6ezxWeU65T5f/+MeRc2rsMwN95m7I8SKG
NoRw6K7v1GtLgtNTps+3BEeC9Ro/00Bu5NTd6uA8VwDxLOiTFVU8sJVWZq2NQ9Bfqae/j+X7dlAp
6+VM8DEwIpo/3kSrhGnMBlYZT3+C2wH8cyCaklfb0gwkvaoJVgXVHMifrmi2bGxoWvdjKqYMW2/p
V4kc2BLadwOYEdpEZ/S+VhaDuq0hdC7vfxGXQ/yIf30ba/4w6Va0kLr66PEBOj/VLFLFQXGKEcCb
AO9KUgrVu5osdnEVbOOQAUiICOIOqpglH0RYRM/rc2kEdKbJVLibSrcOIy4aGg7RrcFVdpneo+N1
3FE2KlKfuegxnHupf73DAfxYaWH0PvGxtu/W/HnyWQUiwVKKLkAIH7OfdSG7q6jCFBHFayvs3Fat
GlzO1iEDYJV5EGzzcBWTecHfsCi6c00+pGHhHqechEPGLIjvEAdVbuv0olPph3DoOyPW1puGmBVH
jnJCF5hM/RG4WeuPgio8IBQipPUnCvB72q5LoAcDkcPA1wIykwmt7q/MuMSQO2OsaRsceKT5ta7i
oxpAzyWNdrdfhsHvC+aog92sb5u4TKAQr4VY0yG+dH0Tl5SQoHRqIQ7ELqAPQYnxiqPfWazJkaSn
NpwhBF7T3NO8EU+wWXcHRCTJJu+jQn87ruZAYZHjtd/p068ECVJdLCjBuTrAqScZgcdo6EfJ1bLH
w8rb3HmDLvGNn9qTzQQV9/NHbEs3EFz+q1a41zM7s0coVqpblEON/Y9Mdz7eAW9v6GfIBNUYfIUD
F1g+PZBvkaanTxyRF6bZm+6IdHdiOxHZ1zLQBJgAJWl2qXC7jPwhoXPnSiPVit8swboMW2ks/i28
i8hPEgcOLrflRMzor9hBqVBKcPaQovmed+DcrYYTkhTInhf6gsiSIj9AkKYWAy9as0frtKe+leu9
+RKaDykeNkgSPkljHV3E5kytZvb48U13sxj3Bl0itZLjQv59o3Pr3Lq82idVI4AmqT98UV4V/5KB
lKykavq33OvRZ4hZOhkQYjiwdriFLpjMfabEcnjhp7JUjoV9nmVEcMC/BjW1t8JoLrL1ujRZCe4I
JyFR2nKfVCn8r2c3RNQSmYcUUwGPqKa+KOjixl/eoUZ4rlqr8TiHu0AsMrpegY6IEMCLJIspl7A1
CY2X6196P/0JAjK2KI2XQE59G+FDc/Pb7svBYwwiR8NYgDUK5nNW4GDQJ0n7YRexRAcjxioCY2kU
9KbP9U9LPSJEbBy77SESPLpvgUEm7wFE8IzdIZK4A28xeKwqihqFcTA4GB1GzHS8qyxx32C0g2u0
eqntSRrUkBJyOfrKMKKKr/uHUSD6OLrTjlaD3Jguh8MKDzLw0f2YpqF5oQqNRfC8uUtwvvZkYxy1
YTLnbZ09WuGcY+ZwNI8SAdqe4XE8Y278lQVpi4o/m/qcXM2KAys9BwdXXNUWnkGnMOgVps1uXs47
gX1x3W2tSx4cXcUDPX5FO0fJUSURxk/kH0j72BMpEC1Fuapfr9+bJS5ev1gQAcTZFF6gbiCikWPx
w3ChsyObr3EfKi2Q/Tc9C+utuNQHGf4sSQ/ExNLh0PM1RKiWcCvCSLwZRbe1KnEQVlHKKObXXvqj
suYjWqKzQum/lnQ6+pWE1JF6EpE/HXogmF3d9DWTvZ/oNyrRZvhpUTIZIE/jux62vkV1C8PKPE5k
fbZsamMpLnMtx2c4sV/pPU9EtlNLZomX1CxFttily6kAn2PKEV3TgPqgQZ0dfgQNc2KdP4Ke9bhq
vg8FXCkBrGy42bHJf773rwV4TB/tJMMfSf8WMpvKcKPzz559CPak6OiTaTQooxyrbAX24NAseaYU
qWy12UoLZ1cNNg9Roiop1Ac9697Jhhu9ts6LidTIze7V1hiD8ewyxPckMJDhcgibs6ZUbxB8z96A
y7unw5UbsK1H6SVyM9jrzV339MYqSYi7QPyecoFAAmoyQM+xz4OjZJnO+07/Vxg2i8o2HH8VXWVj
egmn51casMi6weI4IxundM8UswtvWSjEQe/YEtb2zaIlw6LJvchEhxdyR4jT4YXxA2ieK7iccAT+
py1DXf0jziw6toc2LkEptIr/qi7/y5Ghy6Spj09N4vbXgEQNrlhEawb/hkXDzbDFKveXvMLHU1n+
1W+UW6RAdZPrA+7ULLIZh5hotZPqmUH1uAqJCgTrJqzBCmSdXB2c7oZbShcGvJR1RoMztb0rfOV8
EGi5599suU137F9svlKjpdP+3omKa5UmqGEJhu9THtd4aHVlxDjb8ImMol1JnG15dl6hf4X4jR45
VxqNEPySIjjq89uB4FKAzItmfgFFip5skhkgwc2YZE4NZnR1SMPDByH+xGBysEfefVkRn3yD9hAq
U4A1EuVOF4yihGlkwpCWjboeVxIv1+fqWsi5G9VgnDDItdKCr+1T31xp2q5WEGhHXRY7KpwHoX+l
c4VQ4cLyK+ffcS52gE4clKUqMj49rgeEU4qUSg1WiF+W9Ez4A52pBUvku1z+PHCXlxvcid6fgCNL
7BFnIyWZPBWmEDilYuw0iNeABxVsvWH0VVOXZUHtewPm/5fpKG6aTq90VMCRudOVHjRkqwi4PGSz
XzhP0eVZjuUtW7uzmYCSgee2nyy1HBJ0lqPrzVAqX2BGDzgzaT+3BLPIjsbNZq1q2Jzrd1UJPlRz
HVZCtEYW04uSkwHwgY/w6gFVPjR0feZrvnFuqSMSeJzlr+E8Crq6OB8PlpWy1yCRKXuCGMk8mAP2
wr/u/PEcTQ29oRMw5ual6NhwMKu2Y8yiAvet4GBI8P065QPCvhKzgFlYKfI3uRkzCPNzc72HguK3
6hNToguBGaT2C8DPS54nBB/WlQpHCHsBgrWSWoZoxaoJuE9DHZ/MKuqNFKx1wOZ6x+AFGvrPVxW6
LThrWHi/u3p7FlpEcInbBLAgWAityJmyvbAAgacsppINrLb4ewcBLfORQ9Jtw6JaNE0RIjPOaeLM
GJftfrFD4+HxtuTZybeWefJMsnzbHuELFeutVzHqVxx6fnwQ1tWbdWsRgam1gKMUyUg1FE3tybmq
Tk2eLdrLCLQssbMf8xUTmzA6YVhLrHIe32mXa/10cz9wotNWlQ/+D9pX2E4abDausAlC8cGEruX1
wquJyh3+CsvEyJzty9iSGRFuJ5zChMgT4aMAy9sn174Brx659Aopvk7BQ0VuOQBq3AVbOy/77jGR
kGbED0Q3PekmAGIE20xESRXTMPDBlMG+MwWyElh4f1B8QJk7KfTOlH2lpecboYWcOShQH+V9aq7D
tT9Om6JnkYnpgOApUbHxB+3GY222sZGkKWgj11FryxzkSmQzrCsipQTueIAOp7Ow0D6iKUK88y0n
A+qBHOexRuPOlUV6TeWEESoiZgbwzdw9lycWZu3WeX0VnoZpJi2NdAqu2jg5LepUHAXYPGlGeTym
yQAIxEZ9/hCFZHH+ydtaJmb5nYNrPQSktrLmsXg82Z7BH3tIjgfksIzpo/ss0dw/F0WMqQ+bJQT+
8NFy0ZfTqKHSDoiy4pWPXPy13ZSAcW0+q+gBfpmL8bs9sWlyNbysi2PPQGHnrl15SHZOKaYH9MK+
n1KEl4ykmkvujurV6YH6Va7TZ4d5aizDRkQAC9evlktvG82fLfTS2/wBKdDL5bmlE35MWgXcrFCU
haEOBgFwvnAZMZdLfd0PW30bOXW1BOjbWA0LsvHh6vJI3c2G4L2bTwW9rnMhAnV4z04ynXCaAQTG
374oq51dPHqfKjmVkQJUJLJe4TYtQS0CDuQHfXP7kbc5AR+ncQ2lGynGPuiXkzdAAkWv4qecwaVc
vfLzIepnMMvE0FTJmke8ewnBNR9PLoLoCKWM+NdVfjlOVK7XbrKCCtPSqqoX1JrqWpQrEegBUMgu
4VL2ahazVROMG8Pjt453CR4I0ikzqpxaDwBqOK66w/V7QdrHovth7jfC/I6C0LTF37i5I6nelg8C
o6+cUf/Vc/WkOgdjqiM0a8HceqkJI+dnDoKHqyBGIj4wY9xCRCwDW5I1ZmJ5PQo35CfLNx4HGv3t
JBJHcNitZGOuSA+g/uAgijmAupx3AVYvvHF4XXIL8sYmeXM2Ur8EcAePLkJXobxZPwUzSx3sJHSn
5NtI0MW02c6kjf/v/90bck4itIOKKvPgT+ZjIYOGj3spDKBHuOmevPW5qYZf6810jrYZF9r0fZCD
b4abhIucN3D6YPMkIM++L6lqHppVu6KFhnDJR/U0bd16yNsH0nO/axW2qTa93y4VH4M9byRuXkV2
8NRorApvDagsI+Ol2j086NBpST6+aBzAzRgCjMb0O/8R5+oKksB3N4CvSxaeyWQVnwBWXNqhjzQ6
ktfpatzRz1TPuztY3stAgu8KV+j84B8VAPp+URFmqdUGKfHNHGJlz5pE6T3ku8d97JJR3keQ/4/h
ShCCvq0lin+21Il+grVLHeOflZmJ01uuZn+fWhrLdaQno9L6EoA31yVdolBbMd2ja137tDKjif7T
67F3/8CDwVnah61K85yBVsteDeowxv4w/T/xDJFJ4atutBsJu/pF8zxOVuNJgz9NiaIyGrtZ4ECu
QhvMNjFK1tU+td0klHcAMFdDNE8boj+6xsveVf+34Ei67kIyQNa7f/KWxwTQ0qzSVjsj1OxMydwV
bru7qzLS6dVVjJrWoweZirsZvIb65IPg4RXteqTpuVD1YOZ/hvow3IQbR80gFhQ4SYIfrVG22LvO
eN3wkq+nCs9zacbuUSTNpKR5aHsLVhQn5H1xWpCR5MU/80z5HvGwbw85d1+vnlTA23+DfwNMrP3T
0bS1eHVlBavF2NYsMnR9yt3F5rz9P7JH7m3e03UHyKmnUXTfus/THrMDlTe28SK2GWJ4m7yNz/3u
YssTpT4qL8pwIjg55odNVnh4yyAlkwBUBwfRPJk95lnaKBe+6isTwKxLZ7NotUOmli4kqx8/srmk
znKkuLFcV5jHwDOW1GoQT5w9A+4RkEV5cp3kSuEQFiRWq3qAarteftSTd8coGbJU1mRZSSVWNEOr
we5fn7y0FINpqUxtLpVjhNU2yE4ZsG7k6II31FDOQbpd7KRWHwr87wlfJHTk7Nar5YIomKgw0DQU
gZVPWOhdc3UxMo80S9RFW42MvO5B+KNPMMeeSkN70w4lkAlfmrPgOX+0JDQJy+9fCxbotQUdyD/n
OhzkW3LRzw+0BgthHpce46IBOAZ2SrIPMqF0Dh3ls8ZLasCKPex8uzkiPonVlr7ZbHGEBQsihUDQ
Z2zQSenPytSMG76cOjhCiXuAtSZehgMl8vCmfWI5SaqDoHOj5+LxSCEgRmp7rW+C3GaD3t+NTo8u
SfZ3/eET6nAw1MhKGtTYTU8jKk8y9q98YQFzI6c1PnvdFx1u/bYxMeqgBg0r5WyH/sV2J1ZunVsy
W1JqwvA3I/W6cUseVh7ZQU4ok3flU5TQ5nIDTHMpS+USkLuWp1N2HjA84MBBxX93uDLTz88NEQrV
5APx2UbgM6ZoQHu855rczbgEFAeElP0xgohOrgEBzyLt8EI3kEHHJh6MYkj7Eg+lcwQAYDZdGlPG
55ETug7sVoaYy0LEJsNR2UawdFpljRRs/SgtqxPL+B/UE+g4pFj7iXy0taqS8VHslKjn5x1Eq2ce
9EEl30/retH9NqG3XBDPKqzexGbNwAJ+2FhTTi/N0TuPk0ilJVqE1q4lkiGcZthfyRMvc33viQzT
qwv8L7cIkl58JwXR1WiJYrO40+7n55zCukM5Ih2vry8S8Gp7AwFEKJ3AsM1fEcK3jn7EcF0dq9AZ
Cttu2BboPgAuCLx88bHn7CdGNtAHL1uiSpmhxb1h8SV8Zu8qrErh/vajCUz+Bdf9yTH/khkI7al0
Jmi6biYxZ29AzmQopt7ihb2MrdJDzNFkOnTVGvTPO3xulyoMWAIODQcNGz3WuH2Th2yNdg1ZkQEo
+F+e+xwrVQUq8exfkzHbAkuGztwzhGEWRR38lANSWdDBoxmJZwvVVt7kJswNCRdmTA+5s2p2rLIX
PcN0NTGfZb7Oy3xAJggTWMz4Pnk/TCkNLRJO0jdVCBJuGmg9pHRLiwm23psftxEQoCid23TiSsZI
/P4GXeYx7J31fmb93nKXoFgk3roLxvGsYlQKIchsjm4Jav31muoBt7qAgcKyiAdbYM1Vu9M4EalK
z52ZJ9MUAtdfkNhJlzT9YIHqPEIg0Xx3t2Eq7OrwTy94V6UghlVc1x3bUxVlgf7fAEFvdx0BfMMd
d8WfAqrVKNbekgcRCJOqvKheFPSVbDHnWEXjnSY0ZByEf84sxrmJtpHu7pFal+W95E5luuZy50mb
+OyERJvzkbhYPJYDyMwamSWGlp0H5F8uNggSn6hPUHyvv0qNJexTE1iWXZfSzC0ktFxnA6DmCMqZ
JXtvf/+50y9pASUQdJlN10362YM5M9MyNfBzt8g12TIDJn6lVZur7P8gWOcGXX/rxf6bCPPvF8yv
TPY5x3de5VX7hONRAVDfdEaI3hpHT5+W3IGbykf5pQRbPVWuQHSc8JaLMwFSJG3nKzCLj1DbO6Mh
TWV4K5wyoIS8d+jgLNFz+Cv15/yLZlB1n7FsLMNlsFiISrkd/syhTju8XHT6O0O4MACqFSGTeLFp
SCJS53ZUULaNx7WEyqtgn/Kr8qXrp82i6Ljm96M/VomnBpqoINECBgh999FQujm1i3mN9JwrfEGg
Cu3WpXjbjlB1FTzyYchpG3WmIj8X5fvTiUTJadJalcfQsqUiQTlEH3nur16QIjvus6FKUYVPztyo
oU0AqIKSiNoFQpR/alEUDmPJFNnR1wLFCvIikSHuJBlVD0d75pmduP0Q7mt18GPC6c78QkiMdj32
UsZscRrRUXK+4Qgi1qDCjNNaSU2VdO84ZW8E+hkUzQPIgsnM1GnMKQWNruynEmL2g1/c5hy0oYA+
xY57g4/26hXC2EM9dZdaZ47JWOXVYvJHUHUGWZo9uVLvejXv7qgIJwqDWNOobzzV5NgqaqG+X0KP
hdRXb/7d8zNPQex+4VXwgfYHwBmPQSEhK/sMb2EKeKXdLPmeROIksGwLbcssjqUpWqVdBzwvyEnU
AgVW+NSHMHxWydZg1J/8hnM+ee46Dzic9FMpdNyTrOVE2NN4EZZKysbcPLbpIVKDiTC31f+OtqnP
n0UabSrhA5ip9kO62u/eQvRiYn+pW1bW5xWTMzMjDpqFLhS3dZ17C84Pp4JYG19sJD80Cv2lV7ZI
WSZi26Wv2L3tETIWK9LK3zW4/vTrxJ6KW4gBium6/xEoitIXEbfFbT1kpk3ltz4pPyIDFBiNF13d
sMNG5wadEkDggamYxtsVuQwrmixBLLCJMnZjovOoS1grAH9gb77NBO1FXmurdhwik5yZ6aA3IEWe
8O5wR81a3YR7Jp+Ck4pjOUJQofjwRpHEAlibm94kdQ2CfhddZCcO7ciKxfToCJBzmiHo0C5iWLTQ
0mHpf7+zPOCuEyMzCoReTC7M9ArKwqKMZJAcygiOuBPAYUZG99a5COgrdE6C2PHJ6csISuwUUI1V
R3fWI4rmZkgU+WqyKnSn7ig0PsYvsRtUcTuiPsZ02573DjtHdFfCAxmQ/ifXt8BwGj/2qNjqfIwS
b4/4KHpFJvqofiNjiXWjnIBUNZYCEmH1tIpxykuD2FD4ULMjZIN7OiwP2FsTPPHBGrtpi4GMhCM2
tDpee1xTccWwFnr5bskBOhVNp4hYyu/lHvvPGzG+MLBmumPGN2WUGPdL/EGZxA2SWT4ATgbvZQpb
ZCYyLetDvOXI8zI7JYkGAOH95EdPE8oLaug6TDQKZ86z1sWXOhdBvy0VSXKqqi5A3EeVZ6Y/WjNp
9k4dMxoxTuSdBkRoXkBnlsT0kaShMI0WANIgbuuzlXzyzWW7ZGz5A76vJPqpV/rvF+t/0liuRefg
Cc/sd1cjABEetEQhXDvaeGS0HWoGX4yfVymPjJKQ9hHp73Vhiv7nkgRpQau6p9EaH2BCCObDifM8
BygapZHmVwaqs9GZmLs353XjWgJEF08Q+mvwRsB8PqdeZIgd+8DnjctJQwqhmLjK3CYmWxZhVf8d
otNyLbv2iJnyi5FWHNtLDLnboDrSi3dz6gyohNUaqqHX69BB7AAaVCAo7tXnZJw67LDLbI6tVlQr
4Em+moGSwp3Mi96HeqCA9W9MXK1A8szol8gW6u5THIKEd09U8Nl2e/Uuwxuned/Yeqx3+37LXR5U
0ZVyUd+gWe2DSTMFnr5lC1pmTs1VDXfeB0PgE4+DxQXnUzoSGm2T65LRx7vg36Fozx8FJx8vaRxU
+E7eamhxnGViTBhxNDIjXhFP3OeiwqGcYTMYQ6gbEhWGn9tBrcOijyjraQjg48bLCdA1v865wl1h
X4Bt4MrtqlRagd/wAN3xypzJ4xxkYYk28EvOnj/e3KKN887c3xm5NXvXCUWEk+P+YmtQHm17NSBB
YNzjOTi9CnyPTvSvh7YnxLbBa3npL6yghCikQ8HlMpt+5JUxGec6Navhg62TkwmrFzc5CSXfebJm
wtZema6f0+FuHDD0gQwKLgBqlWrHxUozuIhaPHnuod1/tNWNfCShY54YAXFnDu8CyDmqvAvuuSMI
y0ww7Bst8NEzI8pMwsS4CVhK3bEXjmjAvVUAU5ZVnlCh45eyOY8TcMJAR25YOyQm8NVcIAXsgtp+
MV0Td3DrvT86OAX7fOLUmeZaKNRfm/jJ4BQvudTy86v8GUPrCEDr5+mqG7PSdBqimqxfDVN+v5Qt
udRDKbceutPviCrklHd7TS2OV6ZzePrv3oY9JFp2UbAKdDoiU+CfK/UmTbH7RbskPai8LyLXzO6o
oNrBT60GuQcCl3GwJz9X2p8HpQpakqv3Av+oo5BclR0ImUfMnPCAMt5wjNWAlG2zWik6Q0SMks6z
dAmeg/l5nO4i1UDjS8aTaSpHMyzaUt4hOLGUU/G17wr87g6oQcUw7Kh8aP6jq+dhYA2vR/OHtr6v
GzV5EdSx19ZLDh0WZDAr5dEPvF8ouTuqFh/zc4P5r2EwBkOKHqfASP53ne+G2/TNCaVtGIER4Ptx
WDi6Uf2DHMjSi5QSnBlgc+Meq4LsBiyln0Se5H9wSWmPonEQeDBWHh/7tjeRBBeHpmALGzBYRrsO
Mg/Is/b4Azgl9yzDwexRe4uXAfPObPC8TbjxO3yKLSfjQMO4rkSwMz/Srf66O7kttU6UqnY+7nJv
DlPKu0Iy/yRitRMPJqcSHl4XhI06FnkHffUy/HA+rPtU9usDfI2X4wp208Wd3V7CeMaaXdyPvQr1
Vvpy4gcaEzzh9lUtR5bSFeHqcocnzcciI3wrGxO8mbL4QqA5664+NjRNXYxjIcZKTnzn/uXvy9Y4
x1wg2eIIQplKKm6P+9FJb9ytiK/IEZCjXd6bSIGAvyENMVXFN0wZwaZWEkUxMG1n7GP6zuqdfNGa
/SDHdWmBu552H8vIdVZXZYRPMAeCjH6jyzU5P3EK1ll5PIxoK3+oGdGeZrhJbRPakE7HoCalxTL+
tu6KJARa1ugnV5vW7BiwCEY7bMgowTyjX8CPIuW6z5WUTmyTJNWCQq5OsR2WPrwbajWmhx6mX2Le
RdWR3HoM8Ds+xHNzmgjkqBugLrQaRbA/MwEMrCsCZ9G402FEK5C8pJ9yEM+hAeiBUInYhvyNgpv0
L3BK04BOM/nevcBxfHLLDCN7Xf7qQB+ocKBVXnzUHqOyiQzi5oaRj9jA2/xuJZwlGu0UtOkW22Ew
iA8UINceAl2skb3u79/YaL0Uj1nGfxFj9bsVUsMJYMunLHo2mKI1KYU12CaGyfCptDmmGBC7l5ZI
bvz3Ux9XadY/gnxJ4K+wRBkGJ9wj9VZjctcZW3SCGJlbK1c3pfu32PN00op71CM1okawuz46RoVo
5mqjDJI6U1fVFn6lt33t3HWR1LH2AjYc09Ym983WKsDJhP5Qj+U3FKIhFoDAbsGobBkfke2Ipsb/
dNgrR7Cj4s4vDOducIkzzeHN6mV0KU2BtFycl84OGPy51x8oJnz//7DNLd39pwoXedqFLK7rLpYI
WXCsbZhJOQJyWJN5hJMtfOaiy/Z/ZHrhEDKvByIq7M74JzXA30Z9AObIe7CxNl1QLZP4CxZP6o6I
fuolRNyJR03kOxQDrRR6K069U0zcJOZK1e/4mrXjJoj8YNgY+KfazOLsk59pyvhQlCtU8FZvLbZb
QM8d72or/ysQqPSpjIyKoyNRcQpUjgc7AxiNITY/aPZJBDLNJOmSqtULtxX7Ytnw5d19m6khm3ZK
o2Cc07+MsDjaA4CzLMtpmdxK9EzFhAezK7EELBONtz8JtHQFI/EMK14UIMLTZpQL7Qmn2imqRFLB
MHAKcwGbbfNADlbv75DU9uwWLZ8WHmLhwKNbIAhTm5VbWbihL9F66CN1SQhVsNc87n1OQpAjIBvn
dyj0jOUPnKMuElUv5oXJhBZGf96vreVo7XXB0q2uPQrIcZ+jh/3QiSUD/jMpkEZs1Lx5EyuWcvk7
fGauTxFCVm/aAFLc6fksmtOFxwVusvQskCdRkvTicssLvaHs5HYP13c18IWzZEQRZbqXIQlVqFdV
GLaUJETKGLjSvUI/iDK56+7nLNFHZ0qNJYSHBEjtaybc9cmozpeZJltXvWZAxz27jZ7tJWNlTV6s
y0Y67xy5favFrJKIW4xqkYZ7UfCZbViyW7L0oASgWVvzoGJAg4lEPdeETW3NuojAR8wsvRgu13V/
yiSVyLQqLA/QtoCttmiPWc4uQ+fOeaXyfJcy+c3XrUMeU0s4iYgh1Elioq9/+1+lj/BJJgDdTb4s
3ftxSbQyOAiXn5ChepbidJOOC14plbeRXrx22GVrcONxPrHTT40htVvlO04jbmwyJE0bIia7EJBE
NSwP58XFLIuk0HJLrrCSY2Wi9yl9dw2ZkNyMMD80+EWnJ6ftnrremVcMu7txZppyfkLRC6HH0O9O
z6P8hfU36tIEsPU/xIDbWbPB0JZXQ0gnKzTiraDnxGrrAWrBXOzMvusm+tMgB/4YVI9YxlcSD0L8
4RilTCXM1EGFU5Y5MSzJLC6nFYPjUykL/toT9zKW3C0zx4xBM/e5mga1EgzVV+J24PUeSjxGHjji
5AJoAoecFUWzBvB/G6VVpib39KprjA8mnIrGTKfP2ByCzcjlAzloPEeotultDWWVoh3+S7ag+YQN
eEQMq0f6Ku8EDUnh4DZA6Jfw9iMLeJU1wNGN5fRy4mOX8u0TRvVnILQTuP2XbnxaMlW8dPnLo5HR
b1RrRW+RnlLGLa9A0b8bDa/oJVW0ZKQCbell/FZAQxWTbmXQila3HBxx+t/Xk/E8x23huOfSDmGQ
FJ0Tm9Eq2IemzLe48GS/nsbqyC4x8irasHPZfawgLhTzO7CfknxXglImDX7VQjQka5afSxYzGQ1i
1DhzvPocHz/3Sy/ipNFOcsnfqJKpSCdK2rn8ztPyCOT8HJsh89F6XzcQmp5XwGTkH5aFKuGVq3WD
mp7bhg0SHFtcIUy21+WoyDAvsmcHqBliLisgEeYIo8yzsAN8m0MmhWl7hvPT5t4Ee+WoXPFT4CTs
LHXkph6Kthnwq76KVqa388l2WXuVCR+L8bIagBhhmiv2j0EHcXmrAlRThqMx0zzujh/JqprqpRGG
DxOSXALFP9JqrzRu52Se/F11IJUZIHIXh60u9591a19rOOcd44V2D8Rn1/zLa6avAXQYHiXAY0jC
RU18icEgFQeJ/aO4v82UG8JIyXhIv9WxIceVQoIFasLUc5s8zSdnnupBRVdmw9f38oh4Z7gAG+XU
2JqetjDosko+btSzFozyAs7y1Too7MCodjlX7TmxsfOwkqXcJZEmpdnC2BqTLWpiRoO4nSIhIf/q
YeHavaT/m5/tIy6G70uWl5Sh/EK+oGPHi241GIC0rMbG8QHuoc6XvQELBacjeGqbt1qMoXhXPXWa
N89QNN1CgRKQKwNybHzXLG2RBFoAPJIpARNRoKK+EszzqQTho1Klef+0IGOfef5a5xeCD9ciVBDo
Wktdr0GDk+uKP1clYvueKuAGveRad9K59NYqRBj9CNoumNuPcy2nEBcLwZr/ac966sw0W7G8xJvI
mXFLzzz1GrptRi77pPqitaeTO9R1DdEyT4v7O8eLPRvv0Sev5LGyG1PEw55U4qKP0v0mXs1BC+V3
d+VQKaPhCA+m9dl1IwWqVVuomn8t2YQfGunUmiVtUuSH27WZTz+c4/j/9WS9mzCsymINw+YXxze1
SxWdebk4mYHkMVLts+hWPkZAhfHAb7Dc2OSWrmkb5CfZM92vljPSd7YG21zCRcGpYNur0re3HsuW
TTBonfu7h4o4iuSEA/40/K6Fn/FaHEeieXxe4L74x5nhHILBJgg1KMYWqyS9nRA59Kspoqk2aA8K
qdOICgqCVQkXn35t4w9hSZc8xNgEOs0U5Uuy7muHIazd5QqM0QVtv85NSQcO4ZASwOGc/cFMLo5N
3u841oCGvbds+MXhdJFqkmjTlusoiDimU4/M+1jdJAMPuOKiif/TlzV/5iw/2pxiCSBPzWG3YV1+
KLa4uoJ4A6EKv1LM7otzHAuO5nDHAGEs0mwC8qiIOLpMkHUBpEeg976BGR1LQRRuMFsgmYhFViQr
jTSKGY5QC/BT2B1zZgB0qP/exmgrYm0CVQE3tDSVHKGfXy5kWVts8jYdejMEbmVpU6BKN/wRopdb
ie1tQq/XudQdaumh68is0qLz5ZrWciKh8AgnfHzQ5CWTjx31C86sinsXN/uI91+PCREnmJqJUr9i
2LWuDhOEc0TXP88Guc474Xo1FYN40SXoyzOAYMUPMGTjyXnvF8JCwqGHGGDaAKZ4wrxMMoFCcVng
wFGqNVu3rVeziS1ia9JuUWpJbBVLHfLjks1QnVjzSVLVHpaoi54/4YiaJxYCi6E35cr0iUXNKRlD
rCUofZBVUoiCl63Op7VwKW/LiUTaMDKPJDxHGiGZuo8XuLFdvhLbM3mMLAY76AEnhwGwORtNU03R
M7ToFYmnq8KXR8v1lx5haBpNc3Gw6Dg26JvOdNDCCGQ4q4WCuueL+vQgWmgFstYguqeQAxxTQPkq
XuqYp2j+YioIMhQQH7ZtNLRKf5ttj8Cov6OPb33qGq5dth7MbgLnXQfuNkJIreL8axY8/YucAOVh
e8RN1DL+EfeG3SJTLBkvhdWV2NNvS12AegflghIW37F3uTcw0Gszzn4+K+s5CtK2nWlTt1deNSqo
w/kqRjD6t9O6rmRux4xATHAt/GOWcipjPOkQutRiLoLezYJpuX5KcO+GvN33gJSbaSClKjNgJUg7
ILm24stVV6bMuW2pq1Co3LwGpreeQyicPBBibBhBy6Bs8Y9Y80r2BSxURiXLQSj+50yr3c6h8omd
90HfqGEIRU1TFjZqqFbnCB4jjGt4dVL64c63xqBlgL/AYYZ0HwturQKf8YnUtw6hiz7JcVZUvoqY
T8IbrLFgaraeJ0Ouo1WlQ4+33b/saGwgQ/6WdokHDNF0fwi/yjCUJZeGTB1f6Y35oySmA6PgEerE
/5Z0ufU1THfQ5jnDWV6pOaLwOm59NRuKzcFzpNKY7h2XBDERLUDBrbR82VlYI3YD9s7W6Ox4cxW2
azXPLGjatBZ9BffUvyhOty1CALqcr6lBi3xzULvLnGFiTOlKkxnvzUiIBD2oZnew9l1be2bsjFbm
xpP8COofxg7dCqzfCHqsjXZcLfeBY+dTvHE+SjtTW/ZH4Oisa2LgFhI1e6HIc7ayel0Ba8jkwGSu
DyNv7w2cKEE4/CH3NjNEJzXiYga7SUOttWEX2Pk8jfi2HYmKX/WHUOZu2xRRDQsBwij1wwKwLoGv
YETDgrA6yqYpq4hA/Sd+VAFV6JhN5PGKs7N947Qw/r/MsTzIUdyJRNL4lrznjBy2aF053GNQSjGY
CwNPHEIEkxYgpxS0nNG0bj51GuoYjtq52NzMPxFBtriERMo+AipfvLubbps+V0oIf4kMhl8idktA
+1/wKoDUmLq2NwBBNbKQ+PV9GH1wTBChOCTdA4+dKmpUUYwYi5ZMlojMKVYMlg0znGjKmRA3q9Dr
3K8GUz+InaHmntQOtyCKJGEyn3WI88nzY3VMOTbDtFqPFej9MYf6bK074ycdwo9sjyio6CD3dRar
VFx0o9FYPBhy4IwnGDoDJi2JxOzwI47Emz5TkKnbB0TOCJiwIcJwqVjSD70Ejq4Gj1fNSfyYlfnX
RJEOMLqQ432/SrT3owmjx+WDggudyTafSrWrv2I1ytzE7JXeh0IRuYOSIA4uTcvG1m3O7JoJ4N9i
iHFShfkWbDGMyZhgvrIOgt8CHRKNLwYpoUTJHBSZRM5U32cnCFAEHhW/21cpmN0HU2qYpwrX4HWB
F3XwblsucZupvthDTVmf8RBwcVN7ytlv0NdrX7lTZo4zqzRXe4v50fRKxNlUZwOeYtL9lMWOiqn9
9uTaYAyKyh2WeUDwv4z8GNA9th7x7CaFwKGrPvnftk6OETLtn9bJzM+akq7IBYw35D13qc9+1dh2
WgOknGRYLe4GasKgyJ/pJfsB9YEtVOr1uSNZIMoAsRFTDVDuGQ3xphpPMMsuSFFL9kFGk4kB2n5b
3U/8/jNujzPBcIh7W3vlBxJUubpBrOJL1QXlhmO1mrCOmbgSZJ4+UV5ND1fjwaVS+9Yh3WM0sjmg
l9WAbDCy/FjE7mbK9gsCt/2s4eLtm1jXqlPurdKAGS0hlgdvMGDsGaLVcSoGbd6tQKpIpYtvFwUr
sFfAy+LVWSX9HnSsZgRKFNe35DGcfw4ltlk49tgGRN7ZnJeDQp1wfojoQn7kYc0Dh4lIY6G2ZgIE
xPLG6sI4rRcV0SCYYGHVQlldi7kwy29AflO7mEfvKPLR/GJpL6V/LC846JztVmC0dXnKjrT3CCVD
Eb2/6eXMGUJ9MiNpkQNvt24zaY9iGnKSbd2Q634g25bVDIhcVKEIwPMlhj0eqnDsaE3LHqBfov0q
6xdcU0VUhxIH7aaw98dG/BqLZXUD4kkWOn+2p0cNJfCFpec8DR8FbNZuvZba13hNBhOaCD5zGGdr
TGZNOLAMkF77J9yL3ba4FOQFfXeljY2IRwmFvZzya4Q0sUASz8Akg+SHEZvo7WSkY2Ij4cjx2/8L
B88vbcf7M0YAtZ1H1zZSTtSVjVfy6y35eVaxwkMkr60aytDQk1102mkfDPO9qRoCb1HPU0Dr1POX
DDaZMH1KYn7GACPmFwAb+qMoi4hSy6Y+VSHp9MsJeTireB2qPvKOFqYt1pgTrKLQ3LyBy3/LDvm+
MYF0YsX9XUiXWMEN5M9QpfOVhKYynd/SO9oWXVBTFTG6X+mkxBGsfCThWTzTP1jc4IiE3OZ58BVY
y8rMBC5nxmO0ozuEsgLcHaS3ZXD9daZLWaBA5soJVOAwCpI6AqL7MvmnG+qoUE2qPOF0C+gCTvmm
Bm2fk2pc6Et8kjs8bEbvLlW9/n3/Uagt/zPVIyfPaizsE9XZLryj0IYQMpWbo6cnn3HEKXZHDrc9
VVAG4MBB3Fbmax07HctNM0TGIUrDXpe34LGHHpRp5KKY8z0OqSBVeZt4Vjj+UVrx8EeHByPczwVK
XSJQkn4y7B1EW380uLb6iJRi/fAzvY+C/0qcTZnlKC7oRb26MwYs+aoACQ3OIVyl9uIUS50n2gpV
uxnNkG5pVcXem5uG72PaeS9hyCqWNwjidA3YS//wb8CBqP2FIW2mDaENTs0jRAOd0SA3/kRqnDoY
nHisRA6UCnhFeb2kyeCK/6oE7UXfHYFb80x5UTd9KW1A9gGSfvCjuf8ENLdT/OEgFmgi2ciNYm/F
IrOB5qdZ8tmy1jhSvaKWK8hXy9e5QeeX8u0Xy+B2QlXfkPikXQCDdl5eVXSoH6CEMByw+XJi2aC6
QF971czqDa4B8/JoDXGYp7UjBYxKjIWXkCZ7FJIL0uOoYpy3BNp18/uU0TXpiuwSfMcq3LDC+1YY
Je2r1cxltkpRw5LDzIGLiiTqJMN7bJj0l9DF9wEne20mvay9JZdYwGR2yEU9rxtE+mj8CWv69/vj
fShUgZiWF2fIIclMzigV+QaHbYam072IhayuBhXXy78gpaM4qBdouIWyvYiu+je5QmHaYZWGSmvD
nGa4T5DX8dnecZFpp3vp6OnaNVVX0ELfulasHPOEPy8vm+IAyjZuAgGTYdHJmdTfKdPn3+GZrHCT
oNzAwUqRIoWxk9JTFTAHWqudFAya9CxdwGCS3qB2vIby2tAAT/PAWNOmQD/scnlCI5EGeNYJEX8Y
txbC+S26u+4wKsPZ1hsG+mTu5jkH05BPtUok0IykMmoZudgZDgaERb8ITlcingd06Y1t+KGzW2Nj
zFoxEj47uPFq1Dagau0vVebybLtBO7W9Pv4XAEb3VJPwlAXAEiz/yv037ngF2Upak5QSo4NNyyXG
nfEd5MCGewmVG1btLUmiA9UTb0lTncf3m8fAlD+W2VXTM0OG6bBwzxuZNnP8cLqS1vsYU/nZ1ngb
SqNCShZeN2/b4kTiSF/TTv9ZWpBzvWZYzSarazYdPbCJcwyByKod0+Ox2cP5fMxRcZpw+iGdb159
VYAR0/c6SyMLwYXJ1hS9Y+qgCH3aucRL75wpDS6FE3ttePgjwMsKFFkcfYUtUnv1BTYEyUkGNLzX
WiR+8dqGNTYr+QSfpSYxzagHMYCPFF32Sp7aZ1togqsWeZzjXk7ahtB2XjRCRJJZg/5Ue+zshYUr
ELsbeQgJM4wxNtxmgPUeXipRTqX+FMoVS1wmlPqDV4Rr1k4Ed0cpNGO4bAVHMG2HTCi4Sdwz0sLj
8c37HuH8P1YK7rU+tiU1kz1iihBzpOt2R7gmcQhjipqDW805rhXMwDLpSJEajDI8nHkhXijh1Se2
unwCvPiP2XjEYsZS8k+adV+PSHNvJ7Wc6z7ZVZlde5zHgAq/D25Nkh6dezFpYlxtu0pbPtzf5JQW
pMYQk/U9oRagvKwMmQHaU9odfz0JV0pFbGyX2h7AdD+c45/ZfK1Iw6Ufso1flzxoM7z5LFqm8zJZ
cF78pRMW0jXBRADU+L1fbc0CJXoaEBwffvw49NNLBIOdMq5cPDIZiL2OnUn5qLouQ8r/3jVed+np
N82/rJVaf47veRBuLUq/Gap+mTWq/JrPOJjGpwPEk1tbmzwsSIwrMaI+4DkH9D1eoI/PfQE/qoYl
zO8vDOEsjFpcV/zHyAV+C2VSjpN7b6btWW5smXCTQ09cFnrsiJNlQdmGldb5tS66H1OxB4ZyYL4P
/IJ/NuiPr9O17LjwaLtjrrgl+O7Uie0qHMSa4AXozLpv5zUE8aP50QBfuY4bwepiQ5MOqIj7zpyb
SFd/YckaobXFbbfMBXerZTEhYO2cFVBNTeb0TNoMbtJtqFM5UFZwJ+VEk4tGY2vN6M9bUh2qQYnE
3KShxsVH4qK22rsOKmrEipHrPszuwXfdLHvXXFhnNkEKIlHnlnmi5+7wcxXVIAAB2acUagyN9VPm
tz5GOs1jP3e4hV9bwMjhXHeVrhabbvndITtBxeQy6rpoSBJZJQmGkG2U8u6kSs0riWSS1ohDSHoz
YOHbeatGFzWz7cwwPeNN0lW3GllYgzbstQxskVuw9RDVGa7MEf+XvTwimW1+AvkzIRXBJxRR7JmX
GSeqfNEhxHhLKBNvV5G8547zEtNXKDTwn0I+hoVj7CCFpwWZsW8jTVthBgAJWVbrM94gX9OSGMfL
3bYvybuzrJxuXbS+7QitGXgQPQdD4kRZsPYa+eG7LWgkr4I7A2kkVbQeMitdu/oWFgJX/c1ifew+
vwBEcJmUiS8+exRLUKczpmMi9puAg3bIbtNHjsXus9RHURCwrMNSuf7CR8y00K41Xe4lqsS57zst
BerlmhGb5V45UFCepTdoRwURd/rVKOZUrByKHR/zep0HvNKXacaEBqYdrebiDjrWOiYhT+lHPk1h
e1U5miB5QBT8jiWryDEEbJNpAgYVteeQstAAU/L5fTk1uA7UvITL+NFXqLJV/tw9sfkAw0Blxthm
Hq0yI0vjISqbhEV+46dZ9BP+tXIbNWFycNJMoIFb6r25OBzabJOvkGW6IYj74/b7ULeeBTNie/YT
sYP29PXfdfrnkowIoWHpIGv4fHQ3mSTl/8Tk2ffHseL+m3T0ukMnSiJEAUaDW9QgOgZkljyL3/Cm
z/cC8OnoDadyiX7VB+cTFHB1x4cihVozkBFfjxwcSIIE4LSwEY4ND5HyyWo/EKjcA1e2jcbYabUn
7yL9DxVppIYgpJfazqe6zTw4swwyNNtB2d702jYxj7VtGPBJ2Gl5NILWAEGGUdISFINM2n8x93Pz
KQ7PLFFuMVNOED33bF1HZ8qvKlGhUS/SmMhIoq8CWkVsif38pJu9UsV2f3Dh6ChszDa9I64+aFEP
hsJp4vXWEdvbMcxBwFGqIugDyi/y9RkBtS/YaU21cx6ZIYwrpzdVF5JgdTYc1cTeT2hZYc1UXDnM
QYeHYvkO8DX4en2gdMtyudAhLSLfCryO7XlXfLTxFcE82XODhRBb2fKUhWwVtfiuO5gXDBS1iooH
htDacZl5RDaJyu2XQcdOQqTtQ7iAsW4si73toZ88AtfqyGyeqXFuDbBb/CRZ9WdezsSxuu8MaVgY
W5qxdyvLvrBgKOGZDpazjtGigBrdCK695jjlZanvVQFaA8bQ3Z7dEwjaA5odBQZz21hDnAqMl6FR
ncbUuKFWGBDpRkjfhpG6cVyrdcVY9E3ClSVB47xoNgj7O0x0aO5X366Mc0J+FUwUWknD8Ef6EFhs
IYJrDr/qHwUNBuOeiqgLbaMQAoh1tIRfSQk+kULsY9pBHgjogpcbBUELiyECNkLECMY+6g1VlzAV
yAvWirEeUiBpIQlq1CFDFGBm0Vag2WRCY6frkDSLqKC+KPiXudOOYnBNoO/MF9JHSacvGWZPijIb
bCBYtze2F41/9PX8FSLWpM9FmeaEf7Zd0JNhjQa25FNz1+I/yafF4Uzei5p+pmK6WTi0nehTcUdB
/WD6q2vj/PjkDKhCyxeRrkatVvg3vZdm+e60rqmuTvE7lUgPecRF1yuCejdoH9Rj447x+1Hso0VZ
IgkOtIYcEKlQ8X6ZD0SNzKhyBBZdgQAAg8argdvIoC3M2ZRx57LaWkUWpsGBRpDIN6mBrhnG8vm5
oH5U6gB8dHiJYp85GKUEbhbBIe0N9u4tI1oAo2rraw25rcWN0NsswAn9Fqf3gxz60721bH7q1r6T
ielLV8ce5lGr8QRjXa4cN3rdc/bUsv3qDMKfDzRkbhihLSLhkw25KCYGnJaYUGIRM7R7iIckoOoc
MmfiX1q9vojYoCNa7zzNUMuJgkkDnG8d3eFrrRSdES/HzrqUj4UmRVizA8Ctzw/Tle3hRm/GCn51
HHpbu22ivcByqSlGejCU40I/7FPdVDxhrjojQ7CPznBt1cZwVO9mkB3gfDkvfGGDf1gIpCE8qGcw
RY/hgj1cYAebBdX0nTI4mtBWMy0t4NwSt/vofftKWqcUTRpAMq9o5kCGPOJWAT4fq/T5YIfz8ePD
9/PZP6F56R3A8Yyx0qNoQpsndhBRmnldxzjo1DQbSSQfLPDvSGv7/vUqZkjJtMpP03luwbLBKZBK
JmhwikV9ohDcCnqNdCZnnDVijuh0iixDX0jLETT9rGBQWjdm7bnD1+vNk/+Vk5tleo3nperFaTC/
JmXYBc2qbLE6S1+rFpIZXpSSG3u6klZG9f5tdXYVhW1sYde4sd8We+E8doff6BBTOieUc40hFnns
ijgctLn0WVa/6oZAoCN4+hMCrmDiOCkeY/WT2fd3R5snsVvqAw5rPsqTYbWLdBQ5lFzYjOwRZa6r
OhiggSdUvdLs6G1dMomFVJFU0R3F1zy8/vbWiko3N38jVwyGWePmZEdnTu4DMipViWjQMDyBZweF
sARt9LH7tRMeFbZNownInxSVWGLIMAOpSLuzP7JnkS6JWBSqrtoEIPm/JTF/JADbhNMjjJhRdrZ9
5gXEA0r1AadiaNCZxm5MpXwM0dyRH+Jr1SneyM8wAvlP9I3kR2Lj9lx6sV5SMM+VIOGdvnNL/8cb
sRQVIkeE7alhMFxlAGOM/+CkQMX5KW0zqkOV+K4hAk2Hu3SHjP/ibm2rCbmstz4oL/pkQ7VwCHK7
EOyifrUueIFXvewos8Qci8y278L45cXtEtZefzQYvHB4Orq4WOW8Zmu1OQwQ5FduHyMaP5H5SJN4
cZR5BXxzCVn6LXoBo1rhP9gwWNwqrcG0xa8X0JdvjycwiH2DMfahzPBez5s/vICngGL7Wn8uzu/F
WmSEs3QFJ7TT5ukXbCOjOSm5rzqmKNFqaGkdDCdY68FrYutYBYMtc6vhKjxDH8zYIQWkVY7dcCdq
JqyLnAOQb8vRsrASIKT61OGe27A/na7bWK2lhsA707p+clAVFmwpEHeRy190vxVP6Ho2scm0X0fn
BstkkrNdFEw+iPq8bd+svrMb9NwDl8Ay+e0+yl42VMZ2KTO3mrECWf1eIZ1evHL15FN7GWekWLKW
AOc9cjTTzvITpgOt4XQeWezYUOFtGIGI69EoBFIkS1OtV3MQ2y6yWIsZ8Y9AeJkW7ddmfTfs+uBx
zGljWunSxnZbzwDc+difZ6X+Tm1F23s4jQT3jo7pQdsFSn7KLhbMfGvfD0Kdq4uj8QmP5UOF19JD
36DiAmeZ0ulIWMzErkACwzFvZOrnVD8KMFpZduoFzgl30TjxJ+uKJ3uuCjR3obhWHiTrOYldb7qg
6/JIl5qJKZZ9yakx6V2DmmRviMuHTxi/4F7DRVO/Uf3Hpp6yuuoSpmH6iVibmLKGRm3hLbkf9sH2
lYbc3h0j8I9C2W+qGNDvlRUeiJ8hl9HCUvFIugAOX4ri+K1z7Ib3vrYStrWRGhE6nG2Go5VyEwa6
dMp+8NgOAlPngFBmh6tiURqB30lhZpk+3z5CGOHZTCCl/CYT6A5c1H286Totwtx3Holuhv6Lyi6K
iUFp4lmFLK0B7YzPvq0HWbcCX6lL1JIEoI8iIyyvxFBF3gGklwTWrbfiHtbG0sq5IYwjT/bkcgCA
7to7wKvAyg5a65/kVpCRYArvrr3KqYcNMBbisZ4aAVcXntfYRKLI5RmKrN376M4pw8+RLGSTIlOt
Ldi17ofTXaURz8Q0teqLbo8A2Yt2vh7s4CO3jSNmZm2NbTXikbK/bgOeNh1fvW+b+bLuwvVshQb1
tEoGiQoJxBYKyIFANqbuAS6w4i30JC8tnFOpqnp5Kt68BYkQccBUUlLPoa9e3i5dwkdFG8bljL2p
5MuaVkUROkE0UDw7gPCtafLDXlfHWqsdvTUSOGk/XZ3thM+MzESonZ0endrYewttlNa/VgOD3RhH
cotR8sPTysGRlU/wfB95olQDmQzCb8NgBtMNH3z8YNmxDeh1hGDMOCWchGFVJU586yjjKDMGUILQ
42oMqfwRQcSLtcUgZVYUnVDkx6Kdl8NagBgxBhpCxhzT4UKTc6Dq92+/KYCFDpzg5VtiL2Aa95k7
sHoURAatOJDzBICdVIRHmLhbvFeBsuiQ6dVhgwosKHfsOGOpxQJM9R5viELV5APxdBhVeDecjrch
zQOOqNXBTNN2dC7Gc7l4cNSgNgcvfFlKMKqzitgTp3u0cWqGexmRf69/64iSsV7NofE68LDPGg3L
Yria+y1ugyBcUXz2K46MOjMVdr343sLyrXGO1x1Xi74UXy3n1MloWTJ57UBIi1qf73at3BlzbEkH
1BIjrLuDT22r3Mh6FFcpD5cYBOqXRUmruxXGFNR8kfDzgC3AimNeiQgqAWqlUvj9AVC4VwvHhUWe
fSt/0MuQ9RLcOayqk4Mv0wv2el0U8ElI4LtOaRo93xo13ipyaulk8p4u6B3WWODy5oX2f4KQvc8z
eIMOw6L5EOlEQSwoK5GL7lhwmL3qO3urQWL4dTICo3NU2ENOO5nAFzD3IhCAeB+d33q0HZaWGajX
Zt+U/jSGRbM76c22GW2XbvsyRFYQInefT0JPADUPyEbG+7K8+bHuN2pyRVggWZjJgfjPmVu9euaN
WGjeNvO1BFjJowvZu9MqxfFwRT9vXVTy/oWbSA7O5H0llHRtKbxLMu20FPlKgiQLKSaT/Qw0+vRg
bEoWEN7abLSCWDms1vuS8fzl7CPK/U7gtm4m9KIcEoUQsAwj6er2EyC+Zn8uFCaNJxQNGAxlvpS8
FlVyYjKQr//FuxcCpECRd5kwsCbIP3ha4AGSLxzU8sWiEosjkydv7gdNeqnmlfSDQb0hR2XSmyUG
Ikq+ytvhzso1shJOTq4CLkR9l4RDPxjNxGejs5+6m3p7snAkVt6k3Gt0UhsBJzo6w3cYHa4Mv9tF
0O/+agt9UQUVEEByjZtBFTJUxJuGkseZlM6ufCl1wnR6wH/WHtHiPz90gyawTi47gS6QtAAgN6hj
wLe8Vf3SMsVl+4WyTjG5yO5UfoQQEPOlW8GXOzt4akOYmk6Y5FDI0ChzlISYa+Lul79QknqTeiQ+
vajAH1k+m/S4ajlXfTwv+y5SBMiBkWo5Ot4y0H+Ee7yZYvK7LyV7LI397zCBPiJhFL+jtkdoEKpm
6+Qy2JCHT33TIyvJgmnCecj9+fAY20eB45xFz7SvP4qFXaKjsJkCl6qosutmUBBfTLVH1dysUYmA
jy7YdRdpbqHJ52dLPXDJxvr4/5Vq5sES9FSAhyFGZbpJowL/kX56V9AeytjKPOW5XPVv2pjapRzg
ysLXYTWcDkOngKi0nqOs+CbDO5FUB1UZeXdiQ4rAmVm+Y/H2Thi/PmjG5wqb02/x1UvYgNE4/94d
8RTKnBrpPVl4HSOcL8WlRe/yTo8G0ROElqjme9+3Vof+RElWc3PX5RB7cijYr6NxDj/Drxogd507
CoWIMrrpvVerjsmwV2fjxh2DR7UoF7PUFxlSsjX4v7jsfdMcnv2ufLZea6WqHLWR4cOgrPfdSHbf
VW1aBB9jfYni0GB3BjQBdjprz/bTw5eHwIqDD2mhwWW5E6iV6dl8U6GEPNcHAjCe7WJkxvyBU/l9
sFPtn5jAsbFBLLZgrtC5iDQ8X9k68/ahUWZoPnkXKw4dkDQ3crflu6Ebnq1eIOXDyMq7Xk/Ixies
bLiQ/QIs0vwK9/lAmmthiCkzKjD1dEFUIwLin8wpDNXucTc7X9AefdSwVJDoCK1F23BQnshPpEap
GCkupGrVzhDA0Daa2LUVhZ1A8TRg1rj9ahxVJGO+jygfetwPdTaVyxWkTAqBPTF9jGwhd+9/jieQ
sVYKJzPj+voJ6DnNaKuYUx9KzOmQQiIYMdSTCQnP56SYn9P3FP7HIfMVX4DL5DsKJLzp0UcYXAi9
swKsQ0n3kyHjOAYY0qj8iVSfodHJimZDcpyQ89FRBJfhlKb+Qtoy609oNGxGc79MN9Clh3qgpfCR
T5ahsnoD2a/PVmXPr4dH7V6otOtUtHqdkGqenUi+iwPtLYi7wUNYSjdaN0sGC3N3HqEUlWW+GF6A
tMroc1VbxExMHWA5H6evOBtoQ/n70VvCchBD4CFhEC3c+nIjuqgouvh6A3ZxiBPBJf3qfqYGu2NL
wNpj3yGoVpsOL5cF9y2PACEYTYGW4ZWHfFvkk/lcb4evam/1PGKoOH8J0MKIjY+SqmfRjBFncWSW
AjSXjo8AicgX1EhyXpnRmUxyuRwaS0Uf9LO9G7wd0ykYYegdEtQQSVYD9m6Z8lH6kylxABb715ZP
aRXSTJmL2fsmYD6xVNnEhzpjIcLfodyvN6pd/YbQEU9UhKXAiBg7s1QL+YWhMQdHr7AS2J4JIfIV
M5qK0ANNWay2TyV3byyoWvaSPlVbfuAvu1+w6XqaxLvNeOfc6zl+6ggHg3FD58N7aT5VHtbw+8aD
/67MfbfxF5ldYiXOdfYDcyvsIQFmOPsBxukOtI6oGmUGsQWqD6jhPXFM2c26JBXEghL70yzbbxq7
EzUW6xTfG2E3UbRgbUmLWPcStZGX2870P0A5V8WYaZ8ZjWmDnodt84qH4GqCBqVR/xkM8YQ3cpv3
pmy7akWycSeug/Dr4tx4W+wK8lp9bNAZ1ZXgoA6rXUgDFouexpA9o4rlq55PP8yVLiADT6DfMn8b
z2BJMlf/gUNQPlzOXWHIqEbF9xBMEcQSH8cRmGi398jmaSvBlX2737pDuYG+SWk0HtE158jhInHs
08NsB7Pq8Gep1EThU7fcl5lQvWgjoi2ECoKVJX+m8znXxpu7QoEg6rzvD1yners4saIw+yqcZ/ou
PVHhLCfH/8m2dFrbhmkCZKvS2C/ScuSINx3uG3UGfnIjWOUKxHHWbINwodSLKUdKj9u+BKL55Qa/
6SkvVGmx1GGa2+4pHTVfYla03ChZi/GAtrJxAxoxLz7pqA6GyhdgPrxDD4qPRXLVWk2k+5vg8ayd
vcFNoeVVSfKpV0pXzIPNX94AYkimLxMCpe+dUUC2NAQqIdB4R1Fsdq2L39eMY5x/N/Mlc0GfhrvU
8XVL7G3UIn+29Kf0XnW6VkhKZiyPhqJeATDhDZTNgFQKsaqcdNxxfins4kuqLdZJx1AqFnCR1Lvh
IEks9VKD/S3vWaeWK+f6O4Ws6C/loRZeqABwUL7Bq6E95XciU71xilnq1IcgvRR5U+2vW3MpTOqB
eW2lt7QQk917IE8azNOgkKOdpmTJjZbXWu61YheSQwcMgqy65V1jSezyqxkFGnqXc9g40uUxJGBG
GeR+JQnia4C+rM7DMkOPZj6TD7rIJhXobkdsXNISr9T5WTDsNDvCt9FsmLCHVxqE5rvMuSpoDTRZ
dnlLSxN2mixHwSiOJ3eNENRU0GTT+6rRveDFSdsWAYdWvTtYYNn1vSLHSz8Z1a1M1ANL4yrute89
C4ahl81lYRL2AgueyUwgzqexv54AHo0L+brNBEqHxS0ZE/DySqPPLhYWTrRql9ntWPUPe13PenuW
8okYsTY/pA2Kgs2cOmSg9tRsCtNS4XgJt4JxMRJlOg+feaHORH16onCRZHsvFNN8rDAYUTO29ayl
Y1G57fzp8tj4znndiLwnAyKQOaXkt0/+iSb8xEY6HSJEJIGT0dASy4qvGH18tp3/gly9rA/qTCLG
iRbN6cHItmc58nZCEUhmZImwUZoVWHTtEPc7BBvQs+fYbQcuNWTgrO+JEG/h88t/U/588dOhkVpn
iax/u7uHYmt8ZQlHZfIr7DVVdNuwpB8WYexM2S3wNBO63BcH0sdBwqkkVDA7bWHKUxs1GAgQyrn4
XMkB+RsGMRuwIZJowyVL0Uh8yLeLB8qwU6lVLBkjp7UXWOzy/Vp8EvKQBA9Q9a/uHoecBRCKPuJX
yOdnwtYmJpYs23LCKPh9drFLriClySkSjPKEsAHuyBAaE9bCWTw1kdPZLAlmza026CRkL8oZG1pJ
umFGFJvCptqU8vWyxo0/sB8k6Z0XvPnEXzh8d3azw3mN/Y2fn8hufamF2FFJww/SQmvh8KEfXNVh
Q/L8/w2kZLeV5RcjwoxuM0V8LiDa1FMGVopboGNkgi7azI0S83b6gSQthpq/F2/ElBehGLC5P1T7
sVKT/VTUc6xe12dc45GOBtfXLgmTKb1r36G/GJroO3WlsTjVmEoXahaT0U8N8MQjgXlHmVApzI0n
FLnCZcXATMToZ8JKkOf0b0TfMjN5xFMbwbluU2oENPIbP+mfqsXWRVBcMUCZzeCtCV+O5GGlVOUf
Pmcg+r0SCYGjyPj/L5n33ayDxJ/VfKQuqwmUdyaucwHzFpgxtG305R56CsUy/dcr8t5fqxeSRMD3
vtzRz1k2VCnUt/fE0QP1H01GFGIDALtZeQcMa007DbdQTx9NP24w8FxUJnOyCH/WSyf36iPF/pod
igZqUzYQ/JwVCL5vnt2Z3LfgcmsdFaAtp/ZhV1ashyprB+9gyncGvOHcILYzFxhOhOtQ/s2g3GiO
RLE8ygHiFFlb1tbKEnt7M/Bd+JnycC8dFyYH4V+VB9FHenL2strwPiQIikn0+Q/QpkTs/+mUvfco
axJuChBsmWuNVmJh7c+HquN9l+ifmpbDXp5xo2vILzaqqin6i/ViWUZ/4eKzTnLJdxbDElWUb48K
FOwboAhTuHtmAaRsSQ5hUktWWVgvJ9ZdblXvoRc7LSGQJhgGapSoJMZEUXKYu6ih+WuChdF2OjzA
ml3kmogLX/EVxiXWEaOwDiTw/prK5SlBpcgCzgJf0eMcqBzSCX3R/U2vqsl0SMKzBX7ZkpXWZvVv
wIuGTMjnABbMZhtbkjPmYff2qZx9rKf7+gHLzHItwuz98u9XiikBIoqv0H1d+FjkDH/sTIw5vNn6
bm0Uw4lyESY9ntwLFLrC4vydzNWOjMS2FLESEsUbucjD8DTDmYi46GrskxUSDwkOHPfXBCLFXXZ1
Ah8LANQpCn1JnaaOm9DSk4QkSPVMoZNR7arwBxLlZn/mKVvMp1ECAHkwz5Nv8J4KGS5ppzuNmTw/
mpT+bTNrFYzaV25wbugYG5er0qVxyUgLdqrydmlDtLwRaa/n9AbYATu8BRMBStk0v/xhqBKwP9Tc
wlJ/2PBKxlcJt7LbAXyIHDS2OPnU48DiwXT3YXC/p5LNfSzHjKrN+YiPALOwd7HB/a3vmjk2KpA6
J8/yGO5I5XLr1RxnM2FXlbnW2GhjdENooDAboVLEvPqhAPdicL5NPcXHMWjmgJHvUJvCRJpdl7YY
1etUp/3Pegf297lCBYgxdvTYzOYdMcQLa+4wLiSqvLinw4KNuXMYglsQ1kB2PUUd1hz1elhYfoKP
dYhgJxPvF/14xtKfidH1dOdFKyR0ScMwrDgh9ayjQOP5w6hz0OeRYo/3lCS9yWSvBwG9bzjZbU5u
aFZ8iBsGo9rW9hYY5Skn9Wio1P0jUq5faahUhczcVUAXIRZO9WiiGbH+CMLaSx3Q5T73DxyWmTUM
wZOBpuqrpaJ8sxrU7vz7tYowDKrbnJg/NsG7Q9TT9lWIN513UDDhuLsQCiiOuYSRJQNDjXBODGUb
y9huEEoBXpgZDuD88CWVUqVbdoK/uUe7hsW25JRU4RiENV9Dv4M9dCcuHr880KDWAFw9d5Dyx8yP
kOtAqJLJdM2asAI6czVhJCtNEYaqZdD8/NCya12tlL3PawPqMWuQ4nd8cU/zo+wGq2c+xnprBw4+
PKC8u42nCF7iAZGRcHGx6kGce89wJojjpdUDqmfUygs8QhRAkv1jd5SdCReGVwLwVAjuVOe3CVRj
dQhfderToCAO+Ww/hkAhARpEJlvGKUmDDn6+L7IvI6avn6OHQojzKoupKZN9wEIL2KHov6G8nTuO
v2dATHjv/V7v7ZaAWk3QyYIRfu8YEVIxBzc75KSjbtGqZOwg1X209NDDL4mfc1DaZda/9SGopVi1
PEtw/sTzxcSFxeMbwtqqGdqUulIjvVMtB9ey4XCP8tcs7cHKX8Llr3caFNhmc9wst2eq0NnIyfRN
NyPaJohEaYGhRTOrQwF2Cws0MevCXlo7RtlQHk2fkBCucm1v9VrJd6548Q714AI28H+qCwgsU2i0
EElnTKpwQpyOYFLU2ol4gmgIYXoxCAG7DfNkgGF+KbM+Jr48Z0XW7e9dY/wo+cyOtPtJk3+NR0cF
UYp6R7y4HQiOa81h/HaEB7gPwgYFO/uEZUhKBe3JbjpiErPEPSvjw39Y2SP1GIpCWLNd9XkWDr4W
Cf1Iuvls4dlHOFbEt0hDDd8Cg4Z55olAGQovMzSZ5/qBG+qukr6z5MPZYRI0/KgeUem+iPijGE9V
hm5xS6hKt1OAPTdSMaieXhIGy5SLntuWPdC1qZCIOQ3pU6vazM+xYU7Qc/MTvii8CtCmrCngF8k0
DorQ1QEyzIgGp7xcmF2LYG4GaT9DkkOOIDvPp8gHudkXkANylyvPuARjpsW9myeF8H6wPVvLcWlX
dnFCkPE+SBWNu34tth2Y9k8UHCSfvEsgpPNV+vVWzBUxvJQIHvB5uelixfFihAzrWKsO10YeQPBY
YcZe2YaItHwAdBhVfslICNW44LO7KhZJcir3Gdqax/ge6XZ7s7FRX8dHZFUex7dvgU5bHcCuydr0
lGFj+Pa8/B+3dkwlymwvvo99wp6ffWooNOZuRTidE02OhF0Dqmausfh9ZT7I6Zrec64pz/G2rIB/
MDZLB3G+3nek55aWKlUxN9OvAbxPaLN3GZDmkqCWdvNXNcpB3Mbo/BfTIeY0bnxMvXjgLK6D/kfL
KB4aL/A6/LWSuH9F92AR6umFWLZ+L5r20OBlGudupMr4zJ1kjsj/UEbr74/wH+fT+2Rc252ffHKY
bRNOglY6L6FmmeX9VKwLRj6mYD1TX6ejMu2oNUzXLGYhajP4Hj/gKDjX0kZ5dt6UjRcL9VxbmqfH
mO4YwwpeG94lZeCviWB+sbTtgvsFRnsVB1G85MmMS05vnM+vm/yrxUuazNi0fLVI/KR8w1aq6EmN
KCAP2pv5ku1VCVYDN5kZoyNTIq6PvGpHJfu3/EYd2Z/baSyEyptc5JrFp//0SozvV3X6Wbdp1P7V
rkBciNBcYArxEbDnOhl1O18q7YryFYLOv9SRDL06151F3xPzLyYFKlev/hogPxKNEd5qWCczocxQ
gsntUFlCg4RtSUo6BsQqEWcArHPgSy/GFnNq0COZdrYV8kt1MkU9HT042Z13zkYCXOjI+T5LF6Fc
Cix+ntyHrWmklvxdLmUsnhfmG0RaAvxv4ofC1/NgTenBTKov+lbT2jYy2FsoFgcK8+Sqsc/xo3Mz
HF07zrWCY3uQxCB7tZ/Vx1KfZ/mlBenx4sddVt2svgUsB7bmrA95myRDxUx55Zp8WQD/5Jx+tn7q
ZWxOGOYaLfePBQEcqKpUt6WqLWNJ3emsrtQK10BQuWBKlZ+QypMvcjUSYq8J/2agn49RW815HNjw
YSGPSvmXrllrLI8DdksVY21rB/8Tw35Q8Gt6vlMGrPe4jY9ARZrUQ4szN28+JzfJzwXkRn/mfbWV
SXyr4M6ExP95Mql8s7Jp/blJM5ySxIlyQ6oUaNcRXSJOU8qwVq0lKpEPOD2kXnPEl7D8Zdf9u2YP
btFp3EV4cyoIy+Se1kg4AK1UeiocV16jzOUzECqhQnbMGeUibiGs6w7Cm9De1KxxLahG2xQg7dJI
XhcVuVoE8IEMNt9JhsVWRzjv5zG3L9Bfr6LKGTnouVUgulOU3uFvjAWezd5cLVqUJHFKyPprzVnJ
BlPK5feR00uTpyWQjd50OAme4WlSu87x0TByRnNuIWnqqVJls2JUxbe3LweqOwBJGy407VhjIYy3
qne+fN8fBt005yQWRsJVCW7CMNfo2olWB47d1FGJpCVDlc4P7sfRIu712CQo7z+5lOMtxOVH3cXu
ldyRiA40iCbNyt4Hncf4x8Dl2DsP26OliBkWQcBZSQzQ+CdRHeYzZ1/qaZggKnGXzHV0W/Bqs1TW
/kSFsJEomDr3evC08TimAN+PksFAqiULK7Y3Edv+SgrLY3rUDArlPfsHhxrPE1WvaSFPg7ijJq2p
UwkW57mEcQ1C/do5yY59WJPFCYNwx5Wp3oDh7rDAzufzEmgZ+sO0CzgWus1oYHUz2kHudNQyL0qs
uZDlA6inNlwbYh7klO8ZNc1TFznxn/uDbWLG7JEbFxXnAT86jbXiSmbCOX2YrpSreHSxPncKrQnA
fUK3V0xbCbVp+zPkI+llWW0m2BsRw2ZiLmHNXrSobpDqF94a7rXdypiMZST13RHh0X2XywqdVkc2
SYofbbYPV4yhDg28tgfsC1Vv/jTfOfyqUo2HKiEjI4siYUjrYosCE2g+p31CJySYE6UGd6WNNm7H
Vd5WJfVKmTCatDOK4kloxHgbU9wu3YFbspEbCvAuEH4U8/Gdx4zNi1NUbEHhc798O5cHs27DcpRc
Fuv2PRwurm2VIfKLu8ussh3PmSt3n7RRHBYqPMTRSxOOsmCiD2FX0nptPUg/6ebRqlB1HaMl3+tC
voIevfipRcgf1vOjn4U+oe/VghCmNl/I0DugULbJ55zyrzYi5VKUuZBBz4uUNhF3glvm1ZFeJB55
wGLVUlnSksGr61kPKMQyNWai9/Y7EGngPLFU9rw+hT7AyrPlAYUn8xSRfo65Hrq6jvIgygUuJypk
5bNo5/Wq+P88soqMf8/z66/MzXZMjTNEsFxK/aRAmjICYqoFT1eWjpSqdEnHMfzdOyMRPZjxkbT8
nEadgqy6dvfWHz/xJvSZyBwSz10Wz86ylfMNufBbBcaduVYKYf23mKUtxsDl5ogWdENpSIEMZ8uD
1LfV62RwQuTCKGxxciV0hdSFGYgm/SwnaHJOfS+fPnsFiuLh0YsNbj9vVNmBWbfkeKi8Q2zCDxXX
nYxJF51vHFkbSKRcNyYzWyYN8Pu8jVPGLLyDs8nUwlxZzO8CTaGnuSqku341e320lSP0ioa2i0l/
UCN3C4yWrztINqc9ZryvH6SXPrYU0fMlOWOwEncNEy4tLCyyDm41t7VnhuB1uF1FRDoqO7E2gwqk
41/4/ZUV+0zY8mi6Y9u/EosRCkw0X0uRdxFU86rxT1C58k680Nj7Bd4qKZdgo2Y/m19Te+bZKoAc
SH4Wk6qAXnV6GwrEI0YaO0nvP5gS74Xs00n3EMhHSICaS9lIYKyJseSiAGZ0g2yrOpswCyzm1JAb
qcxrnxUB/RxLme7hr8Q0RyNI1pUfYZtnaxZfHr1VS/3xexKoFu3ew52XCsa3N7wyFyTKB1Oyp6At
tUMXy7meovEAvxGjAp/2Vk8xQt1BW7pzRTIwu3q4zeLiPceXWV5uqsWv0trPvp58PfhPQkVMCHHW
F+yI9vlVlFNs25NhxSTFM74DMh1jGY+TgyPHceNGInGSIaSs9IsQuadxkaD5ctLz+nbvweOOOmba
+lstDxCvIo6sPI49rUNELhyqXOwOYQHzvJFqI30EI9pl4+qg6nICQ3cDiGqOSKswHjVf7DDEAd+n
XI6vQsrBEYK45cleLmsI2/cFNiG+w6/vDaclk/Qw7MgMwwlwB3tWuRjyXqJp+kgtlO7L5DvIzJii
UVozdMNhiPr96Ufl4qx7AsPCnuwpBN3YxHJwtHvTzLzsLXgIi1Iwr4pzGWOvPWqTFjpy/JFpR8hk
GQuIdfCvUTrQwyaOS0O+9C2Ib7vs+LUyLpWd3+5srEI73MsW33dSnxYvuEKnO2f2QhQFzY/uqgd1
4MuYP0twDzd80fp4t5O8wzWhTO+Hq3KxVQGU/SP5bMI2ilIS0z6lQWLiPcWIbBY+WDt/cHhhkgQ2
/6NLNKFwP7Rt9a+sroLt9nZeZuVGBT/iRgLcWl9d4kDHGGwUQNqw12uNh7zrFMNusdr+SfIPS6+5
kNEr5PMB4HmIxkbnZdxjtAzWwKxiUvHcYwxSDax/UNgdx4t8hqc5aqIHGFCW/Dn79f3wtVKfE/Zb
XtUVbmSf/QRGr9XelE8+P3H2NSUAEBVRdApy8y8oG0FVLLsb8mM7fjkoDPLoxgEYWwE75y+LV3Q7
YQ41dVbu0PQoIWSpdrvxnihcZ3Y4Toqc+PJlnkD2SFY95DH6uKoOdc9uktdHqt4f1HubMhty3MLC
xWN+EHVMCWVRYpt0sls2jTG+vGBo0mNbUJ0v4GsmRjnb6ENh4aPr+JwTK/oeQl+CSpqKRlQxwZnq
VNn4GL0qxsR7b5OKb8iCw2jTHHpu4B44qe84kFFWHiQU4SxYG7UdHnVBK7/caD6jB2CjZKshAM6n
thNeXPqdC/UYNokc72K4DZStUsl7AGrr56mAHwR+g5ilwZKQvNIT9vgpkTeYrMZUOPCtNg6lrj8X
T0f4srGifFZiQEzHjK4TDC6JA8O7TkjWZCHqxfDADLo9j4/iUFNFpkWauT0PMiXp4NhnRyqaUrA4
Xnt70baldMgYNxB4sz36X/OQqH/LepHm5r/HbSzvUTnONAaKI41ryNjQkBHtSOcCjenoUgavF9tp
m0sORln2W3N4P4uI6n55gmVM19hW7DLn1bIbaeVFa8vo549hVORs3f5crg4IeAH21SQo27KGDtC9
JEDXRzphHK+rha3DjLU9uicUyxYupBUS9Q1HtVgyNfSveQYbIyBx4SPxfDu0R9qdYGx2MbB6BcuF
BaYQPxc6sJtnMt1IjKI8O1ljzIrRPdpiMpW/Dz/qvfYf29PQAu3pu9itcHhR+ALfrCObEgHfkgz0
sWpfhi8rmZ6nTcagtub9ltzGXBvooC0cqRINW5vkLWdOs/jt/bmihap7zF2KcKZ14BN51/pA7a1G
VvuTgsl+7demD/c4/e0vVJVrmBv07rKp4Ech6Vie+plTpK9hc8amJwQSW36Mp5dGFgoLNmBOPS96
FOEI1u0o78pVAqmPNvNp4wGA8AkLxx4Mc5Ak64Nsw+y3w6kN9cFlSN9S4Yt6ZJE8YtcuVEbsY8Pd
Y3mIjixrGpzlBrjO/P/3d7ZIEtZUFwNjljSt5yXIYmi4CPw36i4gEcaIKOSgMvjwL9Rcx/W/D0Km
95r0ikatHEXWr910v/yHyN1Rsh0Bn8ncFxHD0CW0bxW5VmFenwaru64uKVIkJJ2Ew64n0H1+HCXv
icICmh6DksnWlkMYRba87cPLaBeTdKXtFsZxgPwn7FcEXY9bp1obHW41periSG24dX/H3EcxwPu+
v80YYCSVaVso9FnmXwrPaYTgj3f16f3VyuOGX2h7Y8lkeH6utrpJRweKULNLYeZfADVq1evsmYVJ
fHpp4fmRfKAsdtB2TQ+D5iRnRaUTApfXUx6zzrUWu9aEEh+e9z7VPF7vtKalo3kNYX+4+ekCA4au
0AoEiwTslaA9Fp9h04k22KSJyatQkNdMMxdFgEZRKljXBJi8YT5Q2O/cAp4SD6VfMl2KUYDOZb5u
fJsj91+WdB3LG97znK8FMOB3RU+ROU4pSCPWxbW7E8HkvLLDqRPqrOO6+3peetk9C4Go7m8JRvfe
GLLUMlFDgNUP1PA45wuYKcR9l5WxfjTqLBUos0KwqjcSe6huAyJezoTyItuVhKcAhzw8Mrf0ozKN
+GygnWU564syrZGPc9OPzmea4wz7ymX6chyJmcbvJxjsqXg4qTCkKwUg5SschaDtSK/ESYL0Q9QC
nWZDtiUU6UgukVZk9jBh6zh8M0YYjmwU1Yw+5ysaOBmDhYXzAthrACEdsetOhrvliYY1zgUz19p2
2UM7Sd1kQOa77oVjIMXZ2UMi9UBB19U3lqs2lqY344TXc6ZN+SefVrkw7c7Y+gOjZtInYH9mNQbS
cDlCS0W38gPjpHPGe0nqC2/IqvewzKbvCl/9abBqJEt6m3hIiurMs4lO42Q6NJBIxGanAF7NUeRw
8cq6SQ/1QnXA3u0hKLaGI0PMc5/u8dnBR89Pbkj8kyQA92/CKF5DqMl95egrm+ZDi8o9gWAyOwqh
diCyriEsn+4uKXTcjxVkGTlqAhvhvNIUAVHsEN3hlI1a26Mf21sfGiISon0LDxDJXDc/h4XMdN9J
xZrzdY7UOxVAglJomBx93/+W0ksE2XemAfeUwmov9+S2aQSiNedC3Ntb44vmwwjE4Gc0sc0+pUn4
dK9MpALuJqP71FOMFvlxjXjIVcjXVelFQyD1b/S6dZ3qdQLADxBgSOm6Pe8eiWLFjc5aWaEPZUx2
9FCfZIcfbpYSHbTygSjgv+VhNXRzGnPruNWY5BOa74dzityMii7d08H+/+7PZ1MNFjrCi0hYN+4p
lck4W3dVhlRcocQf1sBocbQfcj2t75auUAf4ct9+lapdfqNVwxWJwt2ryEY4xlpJQcTBnan1Qnkz
P5TA4Y3vKsVWDtdSKZOkgvyCgC7bBI4FxfDeEO2JV1Pg/ZziryP5SthjRW/sXmfYvLFOi9JHRHWl
vZKecyIPAUl0Tjw76ZO5/EkTlrj2DZHsjExzty4Yq9hkSpA3GN1Cf/2wVp5jJSlbHRSDZrCoBeFo
cRGa++xxzB7L3D3bT/VdTd/SBTyPNSuQGS+pdTBInJaN/c64+cbukGZvIgoiuFwwUlHxpBbge6Nv
enUkC19+MoGRj9thHVMw7q4GdkfVvIFj4v5plZiEUcxp9sDEcHx8pIx4FI4+99kSWxZ/TVzFowEX
5HKvs/zjnVX+u5DGiPdpet8SBD5vPoygE5Ltj+uw+CfhKBMEycm9WQ9f1PAh1tLCp4aPrLUj27z4
IdPdRioYo9glAIYXjekZmiVq657pJVnzBmp+rRqzFxPrFes1R4SyNvUrUQRXae82ElV6ioBqJvnT
fHgFn6lvKDDhwtoZ1T0b7ZU806ZL7loDtoNiw3mVxZdD6OsUznK8hjAKFGH1iSFdGhnXdkRiBY8u
q4lqvTt9o5s7VpB+48vpxA2VMCxWcNxE9Z1WsIwIX7W/SzRxELILJ6NMkoo7RZrCPGHY/nigoUSM
A3YVnHb51uo2vtmAAc5FdcXLILiBNUrYM3v/sOv/nNvUzNx18/l0Nn7WsSN6qsAGSon6KTuPi6Cy
YG6PTpng/pt7CF9jL0Z0NlxHwFmt0bk/nQawzs22sV+nhyTqjMQGEOKaA1VT3wE7Dn81LTnI8PA/
d2+y0uagi6MdxVM6mjqVTDvhUsMSMafdnMh00OGkv72bV83KQhC2nXCycEh0NaaWZ3NlQo11OTuW
Gn73YchqmxXLcEukzWKQUuyuHdVg095xCfthxBbIoTLHYunZXpNzkTYTnsc9sWux3z0rpKnEzq3E
LTTeIKwz1s6HnDr0kRMhWFizRD55A89MwGaiCjlV2Jyn+MEWWROhMJzpU/fF540r48O2T9ld22DC
0p8YV+6KQfOmNgc4GhTYrUnhJUhfWqqfMHm83eYBrKlJB5m05wcVMtd5agLmqUOZnJzUuXiyRTKY
WYFO9vXUHHGJa/HnvbbWpjflF6D8ARhiH1S7/ub5CeevRDw4NmEzuuBn61Yt4ngqMTM5Z6uIRczr
gaOpo5WxGPDWQCRO1OUpSfLW8Jqdxixzn1M8fZeemz7g50DouKIXIaeLcKpPfK7fCGLjJIl2P4D0
GFrNGJIk6V8N0nF8P653/ZzBLA1f0DphU0DQy6iQTb+BNubl6GRlFnixMySe0PZ0fXIHTo4pgzY2
vHtFPw0/X/vQdYd8VaCD3qehqObOD7NHzNWX9jznqF67wYsSd/JipsTOmh9/Y4gheQTXxLGKLaEM
q5/IKDEujU43ALXl6c94IztFWuY6S2+fM7bstuLgTMTAv2dt5qySu5/2g0p7RKnrVf3w0Pv3ENam
FnBEYYm4vUvbEtme71l0dhiOty5q6TTlCnbckOGWvE3XhnfFvkiPifMXgsI8TTeo4N5J6jXjB4Tx
SOgJcxcDy3C2IhG5uWuQOOfmvQZi5QYXY2ywaqdZ6NBjNiXOuuMCXHslz+/PnL93GcIv5Edi5/wn
m1kMS5sW8LVRyYV/o8KhjSwR+uSwrINrhon7FZS2LBP7oPacfRVXDlt1H2XBuBFVKlxzyMrIJQi5
hpslCpg5FRa2s3exHWYcYHI11Sj4n1AfWf8kA4HdaJoV0JC+JS/NhpyYqYqGDJXvYFhWPmaF0Rjv
lxfUzqiuxnC2Qc6c3xBeQHLnrzCrtDjzVaw4TsRaMsWoBx5IUw+GkkfirBxnDS5m89e6MxK/5jmR
7KBkJBG2rSm6rJpgad+aGAZ5Tu2Lgfbh3q4n9vuerxJD1TcPhi82oR4DGxdkO2V8zzNLePCYKll3
MbjW6Xrnbcz4D1oiXABxeMrFHOBo27g2E8gioKuH1YLp37keoz4RRQoX5Jb08DVt4O6N8paPFl+E
xXYuKBI8RmAnDQWGaHnhGRxgnJKfJmHbn38ZRcMVH/HH1too8ecMKH3NoMxvLwR4+ngwhjuWeAqH
zCaNyd3GpvIaEXbdNVBL9dCoUl51mrhdtfhOo6vQs45TmPmKAqVbD0HOVBupSJhKBgCdYsbZi88v
dRccRyncSDZzQA0knhkhwZMK2MMLqcK1e/1/X4nEVCi1Qvm6hPfnvWFsLMLJ4EQF6HEe7CGP3kGp
uvjmIp5N9Rb8nCf/4yUz1NptSzfiKMM607qoiQ1B6bp0sDAn9VvI770sWHctKs2bI5jSuZpfCnEv
y5tNm3dUUTwmP9hCkOnbc49WMd/2780BwRSsPb/qpw/3yI2iLfmaI0oo7blmbOgeaVjxq2qAcsHS
UwTMtdXFq5Uuf7Xj11C6I8M3kqbp1fEcSPs2AIbRBPYkpeoT1/TcXlMJTn3fkj4+puGeJzn5LqM/
/bNuYDgZ6V2Qt50LSgtYQb4OV+Duq5BlNCulpA9g0TOtABve/ItDInCOs2s2vFQ9Mc7QzSeHb5lk
BFPeru2UpRDAtC39hINzmsuA8Pj8VE4n3+iJGsFKCe3xAAPbERx3F0Ak1h5Lhg0iVcKWvP5U9EUi
OVB0WTIzsPTsF0FoQ3v7t5T+i9YGPZ2MXKnWAOnWoaBnm93JYWq26e4xrpR0Xf5ApEYrL1Jmxfim
kcsHx3Pbw5KQ2YylXbQYI2z+HkcfccDF7N3JSfnNtkS92iK7Dx7Waih1ooHxTy2/HVSNzP0M8nus
lYuwEGfgh+R7IIkIsxBgBIuELvaABkOqlglMZo98TijBNEaChByeZs3jShhq+kGaoirITu+WtPJk
Qbh6b5Ou8KeYxmlHrMfsGfE3bvel4vDdV+KNYtNiuHW6jQt+c5b9gipOiiwPPZ/SLe+injl6NWOE
IqpllJPLRRkprHRz/GKSYFHI+gYcB9B5sQ4dd3rSF85CWhYpyWSEF9ZC5uathmU+mFUqY8hxgrYT
6bmadl0i8KOp1XJuRAbpKJZCuPTW7VebmqwOU7rNoxDSUoxqmnigBlhG8XKyAnkcqTFd0u1Y6kCo
NVct21SlwP6P7rQGBS5Nifq9U3Ivh9UFpp3TcG1KBzoaf842Mc4awScMLtaNqnr9QP1MkjX+16Dr
jwC0MzXzjS2DJFX8xJmja5B2aDZRyV7onpMLjbGqf+Gkov3OLiVPTmFRWX42NwKrx1fr6ClYmx8q
2dnOH6LI2S0GydsbpNLKfxKpFZVyMJkuE7ow5RLl+6rndJbrrN+tTHlnzOjQy6to/FlMJlfLQPVQ
kct96btd9Lkm83QuvyiB7e6EREf9WiBqmZtnwsX8Yo2k5KMumpVAs587+m6RMPEOvUqFf4uLP5/B
RHo1a/ZQtTX5/MogzHMGXBPwQumqtC+1NurfBQBuaZOstwc7J+Wrh8jURT8DLPzcaxHyDCN2I+xV
8rVrFbkGfQC9/qbuEGvun2Kt3lsKdKfzmkle+53h89TRlnuQz+u77g0pqCyYI3awGfWGaJYNSopJ
gwthg9prII47oMvUzL53Kd2jqcpEq/YH4kIMHtoU5tXWA+rCw8R4hgDQfQOTXz6cyhVbxIbYe1x5
Q4aomFWRYVbMILckXA2XVrLIVX1E6fRyY7gy6m6copLOfA1SwmPHAznnfQzLTxw2c0664BUMOfID
QwE4oxA7dnvtXXydSLGtfxjid2XVjO4EZrTf7z695r/0FfmmfTOgLN7N2cI+T4V8rQdTNfeMhePW
THD4oD5x/KSyRh/KICBSK4n694xDLuZdldTZfUN3Az2DbAEJy0NfaDeTVkYbXvnyPnIABC/1Az1t
JqezlcpvaTEAWyDvTpSGYvfFMMhWKudi+xyKi1N39LKIaQPUzrzgd1MtnBOnZykR7nmxyQbP7nQQ
G53Xvcni572JldDCxdZk6x7fZdDMhjaY+AuLRdVxh5abAjeG91upQoUPZYx/JhaLkKxEHnAwiRMy
rFYpUEvcA8mCkCgBzIreiVhfeJCPH6V8EfyeBgzyrsTHBa2pajg+bBMtnnu8dNv5yEFdrti9Z6h1
hRj7EvQPQ//n4G/ZvSHHphDStf6MTlKtFdUkHJ01SUwXNU+IzWJhAX61HY1+mQDku8VfB79U3c7l
Iu+3C/aqaA1LxwPoVLzhrg+By2DCSSyxas2fLy6d1aD2qH5k+vezedNKbYfJkkCwr6mMbd9/u+t0
6QTsjBCTM6U1TQyGxlXaMLSl3RuAjHkl/vtb9iFgSpSMrd81T83+O0koPlWl2TiImvZKrOh7S2RA
ikJJ8T9zu/9fj8954QrQflQOtx++dFmgzs/PLyov5FQESE4V94gONcmSqmRmtVrzNnFqIf17ffux
3r8rFORDkBsevDgJXM5xTMPtbridkrLnEkjX4CSJxcxUFvxaNCkgODgYgThcTzrUt4Q0HNBr3MIa
ljiMpNR3IO2sME2ivC4A4fYPi5ah1hE8fk+Aa4fXy5ZOnfE2SVg9s0oFiUKNVyBxIBgDfcez+wNG
Xi2sNz9nTQp+GrCVkGohUclRaCIJd/c8iAGavRcIPTMGNvLmyubD7U/y3AzTD+C2oc6ZaecADw2Y
A5qZGsKF+Wyn0k+9CL3vQC89lreI1GymvHjA6zRAI2DS03ti2rmbkfJ7TnHSlHZHIyVMBCeZIajc
L4jyZdm3uTUGMnB0Zxz9aC8+2d9wzAa28Q6+jXsfMQBEmmuRFY5jYgBzZ6sCD5MXp6STHa96Et+S
WDavedDbKvhnFC2tsyNfTnTBvmwDVwKtQ65yFGF6GIY9xq0vy/HlcRo/aeX7tuvtwKR/z/zUhBYv
EItfZR8Q+7AzvFAJUr9K1lvkpM8SPyaepa3pRGOahfYhmw1Cvn7u90ZUy3iKKdjmSo8cxL951vZN
4aG3I5QExXUHqPPEPZWw+Zpk/H89wOvqZlpMvxBx/bK+5lybuVI3wNNjIudzPhMMMY0eB95vUjQD
bHrncOFqURJezMxP9rnTNXYMg9bRLdN0orA7hDRhF0FvNqRto4hHfans0NvmyfVIlJN1RKV36BqW
aOwZU3ew5jhmQoT/ma5o+zeWvxd6VcVKHur6haZtoJ5StxAl/JRzoYXq9yL8OpRudKIdjRgcYJfd
buzzXx9W1urU2k3EdHPw68/W2NmgcBYwJ9T7qYbY4cryO+8a8Z8xytpTqFNairnJYqN4TvVbQ67b
CI1XDJ+gEEazGnYYuJ7YvEn9bHrURWMJu/ckrQ8uwa+k/ricjqNIVQ3logmxLpflpuB5zSTN/SqX
MaQg2sMTZ7GVeEeeyDAwJ/FKjzuyAFYL9ausNL/albeZp91yNRzzfneeEt4EJnE0hgULrSL1o6qL
3PuKEZzOgIsJct7KrixFwNmnWS6X+SxaldIpkMrDq1SBlXLcsrmF01uZqqhz69me+xYzQd02ex4A
9SxLKgJBXLMAJeV0M3tFRtZBADxjmzczsuYg8wwpgO43DSI4mkfYjbTmnOKvosFy5zBOKPjxSn5J
zQl2YGINc2GRXMFbp9yj0c1596Op4rTg03xjW7PGT2Xtqf6An3xu7gfkso5HWUL/vU/xNVYXq4df
gou1E9K5jqxrTM3XOfSklrJfU5oUm1C5ESr8Ig52IoIp7knRo8ljm/lvD4/mVteu6G20BkJ/SSsg
VQPtkR/NJLscrt1V2yvy9s4jj4aGSevlSkkPKZpDSFkMKxIHw8gaRUNk+ZuxIU4x4MZxFaTMoP5i
xgR+gceG6b9fRngS8bTFVeA044XrtkyanFJF9mR0iDo+Y2apW/q8VL+3Tx7OZ9trfxpvtUMkyeAS
ZBbErgSQ3w49U+bFpoZmmOAl6tBYLLlJaestVE8LiijpdrSNFf54jFZaDSFvImYzDGZ2bnSLkuCI
0rdCTmPth/dWkIoyG9tVyDPURw/f69nH1jKU6YBxen2h0mGFdb8LB00y1Ri+VOKRkd/WfpMTWJEv
W1BMl9TehfakbN7/2liuTwSt8gug0g7pwXySBu2gvR1SXL21x//J9UBY3Wk1rR8fHWQKaBfuJlqc
7b00iYG7F9ZiRumqYR6m7CZQbmhMBYHvizpX4VsAyMnl48mm/eQQSmQQXL4IWARIGjsUiF80SkrN
YHm72N95K+/hUQGmznPB4YIqKhqfFswMX55m6C2q4gET3xu5Z8sqRmrHUbnts7nBy6jFwIVugUad
6C8LGrcEdkPAk/CWvpeXsSMTLuRMr1KtAfTRnm5msKnGUemfWXaRwQQRgIURPqWZvahkrERNBhlG
MWySI80f6ghVMnnFMj1OnhptmK3PTvWbw2Wu4umLho+b7mu9vGgsH5v9dn7QKY+eXeSPV31s3HbM
Eh3EEeSj1r5g7h7wiE4je/IXdhOtrGVD/OZm1dmfPqaGMijlfkVZqFBZxWV9b3gJFXKNr1Iofkyh
QOnkZoDJ1VMx9bP1EMu+Om/GjVHTmCMNxFYCjTU/7I+yXyVZx90FAWetd1YKp4GQvGWJOfo1RAiE
Ru3bEeuUgBEjqE5CAbTE7spzGXKU/GEm7/Bvxe9gWmCoYD9DyDSrcH7LQ9O0jvpteaLk5Ab/8E77
rzgJAaxmpZZZgMPA1aYssRAMUcudlG76qNXvF60G2+yBpWPxIhdbuA+EUxepf7RsgIuK3ZAK1JOH
MOkhG/5WLIQJo85HdIrFZXMqBIFlrBiWf0kUZidxz7qMFHGdkfVjQZfkHAaJM+FmM9tp3qcTvg2v
/bIABMOdU35qSwpkE20muLEdHu93PmRrVPJiUras/yb7Nh/QYOfKRH1dsTqYK1HOsWaCuUl616Gb
T60ybfZAlN4IlcsguNWkKcK3PoRHEPD9oIQIPmMPCPBZQ5Wjl5imWcNOi96d8j6R90YwvCGVtdb3
vVkoEeRKf82PJwKu2t1XdDaUaC01PpgmyJZ2Z5ckcIt8QWen0CNV7NjwQykng6Ot8diM+riqsJpi
OjeLctYfmWzd+CSeaiAD+Wv+XWnXN+jLjKPximF4sH2zaMr5Uyzr2B1PqGs7idnIUoBbWmRFFlq8
7rTxbYW+rpJHIy4OnvYywjy4URuRBNvslE8KkEdEy+S7XfhQqlQ4IBpj729dlsjFtsqigN7XguQo
GPozPtmPEKTX5OVJSZutSeFUSJDnjtJ2RaTsTknKWFgxcn3JKfZe0CUCcSgeqUq2QLQIk/IOQJZL
+xw8xFT1hFXsRJyOUOinqDWYShd1FvEng7NDAKdUhvBYovfWbQ1y7ANbIx2sxq0qAH9UCblUM8DI
pduHf5YKMlFqXEg/HF941Cyddr9n6HtgpF3hsy/L0AfyLIRH3a1phQrNZDU91zBsvkqE29vGRL/G
CNepaqSndbzg29VCI08DN8IxL3x40M+xtb/uMb8LkcxisQ6b+oG9T/BFcNQM1h0JXiceFPPU90BA
Hj3U21hJC4QlNZptfgBbbM5Gccaz+DbGNNWEexv4Pheumjk1UTTERl19YEJ0LqkLgvo2bUeul8KI
+VYWm6ohmjmbni9on4njjfPucUnHCwTBqHZW4BznKxqU9RAmZzsoFUOcDQUB8GJU6T7WBYXAMx60
7xBzm7b91ep68eAe1nTHGcuGqssNGKMeJUB2EMwKR2v1/z1jDvq2EYKSihwKwj3xoB213K68zkNI
w992jTuUal3mvII4TME4h1Uj/Hu1BXOk0wE7rWlincqCBKuqx16WhXWSqcnd55PNQj5nV2tC1IwB
AzpcQ5AsYTnSgbrZbchkgttoWlWhtGz2bYf+tw4HouPkXEfFC1dUi3+nmPkopNMpUPFF5xNTLX1A
7kNjbmyUH89MluZqlk1VYL7mS/edKIAusSa2b2lPD2Z4qowZRO0qO5Q6MKAHgp/2piRYyOwovR7Y
UgaxnpPgsaUZgPLRsAl8Fwa8sPhlHObcACXyDMnQaFcUQBBh00gQkWpvJYmtqziSp3LT3wW5H+p+
KKlyDf1301pyhoDLC1GMI91GRFLRgHSGEsDow71odLKrAYk9MFx/kWwMQM9mhnbiA74XKHJlYfUF
1HHTZmtT96GnUx1H17ekGz7M6mkBDGfEYOVBGIqXH1gb+xJ6Xnn5VtJblzJMDFsv0OLLQzNQpQ8F
xdfIHRwmZi09S65Vw1Yn66dzz+Nii8aLr2BmZSHAUU5UxXoisszd+fdMtoYSCFtBnIKr4Y0iGiZ7
nNhh9oFyQw8zdpruk7FOoLU6szL2yS29raJbrBmhMuMDuw5YB6VbHRJAyjfRpH9mDh7cY+fjgMYb
N1Uj7vfHyig9kUxkfbPb9PvWvhunjmq8AOeThjM3/3E27NpDeYL7SKFCRpoiBrKcAfqufrNmcyDP
WtK6nc3VzNg6TRrye1ETRJZmuLfeRw56xM6NunwCJiNR8eUPI49KVhVPWTT5YXBH5uWkQIVOqFNR
yOlesW93cj5T7wRkqYMG8M+L2s0uNjItbpiv5fS2RnraoQzGPtGzN5czuvAlAPEIcr7xvONnF9sw
zLiMe2Gf2gZUq/OtzHVZ0mpL5NuSHkT4PKO/J6Ns+qhw+flvoiEYL9w/1XSY0Iym9TAMm/h4R7jp
04xwtsa0uF3Dr4PC6bRnXmYHaMuXvDsKvH69YWxaQfpk13OQ9OR2rWYyglgu1H+cdal/1fF9YzvG
94uA38+TqywEpIrvAb9b+srY/W3VpuUpAreZc5wuB2eQkY+Nl+yyJX3h69aG+p2GufePMeuobc8w
IprLHyfkcJAK3YTnxTMXYPs6+DF5kCSJuVbaN63R6WAq2HI+FdgTd7jrGsxa7DIcXvIDAgWkGJv/
FQdN9wc3wN+ffkRDiK1izpZej6iwFgMnY60MGiPodaS1HAaLEDuPvGZy40NVcCVVjw2/tj1I6kzE
Bs8BNeOihEDblngMxg/7o4E0lhGbqDlks+fXpbqbuVK7X1nQv5l5c74qBF4aMXJjSPF/v2+sfQzn
VyDmPPjlTOy+zmYB3Cew2UfiYVAsRwti9XvTDe5B4bLHgS9sQcbdcsxDX6yb7AhvWFzDkD4YjES2
0pLzUUpz4lHysFFOF8bH++lIQLKhcQ1uhj5xSa3ezIoJKxt8vlnYUVLVD9ForMsy/cpkyMe5TLRk
CTzSAZ/SFUW/vQctgTAaYIjSJmi23Pd44D0euYyAzan5jbrLGtMhFHaVJN5XyKU82UamI5EVZ3MD
70TBbQISYpC5cJnXX8Tvh/K99nHJAkLE3G+dfLV1Wxn0NapzvUhKdRVxZTb2gKxk+GO7SkdTDIl3
dkqV7gyfbbEfpXXd8mdpj7bSp2iSPM363WbSylbfZAoL4ZaTdO5cvhScuIb5cRqwvryEgC0IoZyh
cEOlE81xYOurZgMZ4fQ6ttX5GrD7Gt7/ArP6nhMNYBVnsPjnGp+/AuVwJ25u8wLEWtsunAyKLsBh
TvFIqq8fZIcxZw+DUpoGTmztgvemVNXS9NIGJq6PXbNISCvExbPBIwc1L/LOzcxAYF+y20FcFHP+
H+iGhNi/tl7ARDJsfFjIAarYGK3N/QF0xyPvpLlS4x+lVZNjOQIxqH+fw8H5H4jQEH+6Z1r7lyq+
r5CzoTDOm/B2QOtUkF9GPocznRvESbX0x8gVYYfrHhN0PTToEtshUvRFBfOjdojjhDW+hFwAA9IO
ayEbjAjWVbycDlXpHeWrI3SNNlr8jdq+sLC8/S9BHpcvBhVcOZwf4IlPsIIVZlnGd/1LVdXWMHVj
27enpsN5Y9VaYjux6gaf7V7qGueZr5U+RxE8UkXJ7XaS15fL0OzNWDuQ1PlymL4axj+AOs4+/ixi
Zsm/QBHzjdRUXIisSH10xCcr+cEWL9PgitRYtG43/krHUEuSqXi9gLfo3MTJAp+bybKEHh7+vqEb
1QnjkCzpW4HAXdZ93SBw7dj5gORgXaxKTbMRfzIp/k+w3Mehw080qWWWqKYzgTi/l7PChPC8Tav8
lwz+hu5gWLpatlTl8iIi5BNYlOOAXjtVSbJWaQlyT/eBPvb1Mx+TED+p9tU0C85z8iBLeYDaXKWJ
dinFCRCaBYMavN6LKKZbtaJ/8QYkP+rDk6Iqm8100fcz/F5J13RRQYdyD4juOkJZKdXKQ8C51tNX
K1PPtnngMzxFKYl3osdX7ZKt5P5NFq5c0/bz6Fvfv7k7SIZhtcgJKhe47ZHMHUQ40Mr5uZNHSRRD
jfO/FUOZG9beb1skqWAVolfhsZwsKrUeTdCVhk/Cek/nOpp2KeZ331BEePC1R5FyQZvhmdMdXAj7
HRpOALa3ozNfIGNKh36IgN7lnb84khGz3F8tFcOrbSbkf+UStusfV9QY7txAJeJW2iaS1zBhZ0nf
DotFHpRAkTtPvUSrHa8kaw5qzh1O6R0hCd+lTRMHRPdhrX5paG4VT0EJjtlwyoyuJ8HWNtHcH+OH
K//e3K+pTTgrb2lcbeqYRug1K8xz4bRtmr+JeU2m3GS4sfLU8hPGvUf7YpQ8bH9MkiZ2kNpiPM3h
ssasYVFzW70mgOBAyrH78My2wEdCs07b04Jox1hZOjusPYB8S/zA62bu6oWBGRi2bZeIr8f3hNTI
OsfZwfANDCF1tdKuT4D/5b7kfwcdcTS6R/4eFOYmnIF0Pzj9groYB6amW7I86TvRYNRJGtTIDfH1
Qq26DlRW5UIWHmHKczDlDK68Wc6czbgG+O5dICqY22IAs8youW61MF0MJ6tbp59W3ziRurRBNe/M
tAjfi33gh/zFYHh64BCd8hVFAmL799Gz8HuhUEY9tN9VV3Vsl47t7bFbbswWXvpKThoP5grPZ6hq
VvZH/fPGzS7DMjw7DVc7MgcW5f5ujyE0mQB2lh6ROD4QpOXV1fzjWCCViq/Wc+KEh5Ofo5S/CNMA
NoRHVPSRqrFAkccX0iNDWJS9p3GP9j2tXkuolqLGjbB12G0FNnhvTzXlj79CLQitt5nzFKdYNoiU
Upmb+vvncBF9+v83rBTDrKVDGhsmDspUlAavFJDR7eB+GWPS4Dw1gnz53vee8JBID7IJpx8vTMS8
149cszRb7qFGgfK51UPm7haCGSH8XqMIJ9+/sQNrJDJYh3Gs5LvDeNH7jKJ0lqWH/lJU05txpmRC
r2/YKgF5K6VP43uvZe4595Lo/pM398SJc69aVy3rJnphnrJs/VSYrh+B0Oi2eUrxaopSDiBWV/1c
hqkd+FE+4nwnqffwc6SiIlugct0ENOEDcFHjNIOlSISWspNhdUrkI6oXeXbqqjUZXDMikRYBT1Oz
wm6kG1kf/8/MjKw4sCc9adbUkJtr96Nr+VkgBoVr3uEw/Jn6lWaaitQmpJsHbUyOLQJ4xonxYg5K
3KnVUYGNl6r6CxaFw7aqud4hyLa+5TreMzj/dMenEwWEESs7M5zWkcLK84CEcqLUesfHX+ETr9zY
Pd5MhDMnkCfpsIBcsINzuMjtDP1z12u3fUayQCSQYC+CoCJsmd3S4gT7WzfI550+VPFZq3elN8rx
PNTMILAc+W/PQscfx1A8DVeGftFxW92uKB/4iKm1feFE/oekI985/B0xV7mx5SusOIN4ILe+Baxo
b6iiPjYYZSDVKDNXDxBl0Aqlizni0qlOu/BvOLijUJSN1VT/LQ1ilyscg331xJRC51cZL9n9zmVM
Lz+mbHaduuw7djSlt4PRfWgEbMeWl57pVoQ4CvGop+zPBdYQGVEsuGrHUKvd4nPpN5coS8t5ccMn
Ni9e0MJghRFFg8Z3/ULf9OUSlqTPIe73o0d8XgZLUnzO1saX0rtYh4nzmCGzURJm/hKWSX0OoFGl
bew2tt42CZ4NepZxUp/WF77XGk6J9AyAQHBJrMQLcI1DGLuH/w4B99yuLItUX00rpltk2vHkYImK
VcdS/5BG39F/vXMFQBrA3F/MA2lVOQwVNq168K3+uWdXn6xlCgaIGzOC3wl2tmqYaPO+qR+WQjMu
RWcIDDAHrwDeFyF0nRJq+DEBH+qnggXh9DaB1xTG1tikyjI+JAQHRHmqvnsBUQrQpyLrDPd0cMnh
xGwyowT7h/dP2hNjGDwp23tvkgYlvjI2LQTYHl/SAZRtTt5xSc9ZiAEAWyJN5ZkgHB38b0KXCkGF
6IrnvKwuChzZfYELI0/p4d6VW/SS9hNNzrTe+Op6w8bT6dzAOHksNeWcZZgyTMuCGelqX/0B9peN
rKCRPy6rqKN+ZJDSVzC75I6eKYeNUQku5g62Xv0w4TuB5zNxfMtkOBqbpV2TTlFjum3C6/bnf9nX
KRresMW0Gcz3tXOuoyzco8hfjIotFTrelJ79i1gvaHeaUYxBar+AcbkFA/cVVLEq5/rwSnCXT2U1
/2lG9Wp5SNVrMR9sASGWwfBzrSRXZKA9OGET00Jzz1iDgr7f1VKKGyzpD3iOHzngEhsfGMm+YEfG
V1DFRDePrTXUYxypvpiQAyuDKCy3wXvyYGqRNaWB01SrVTEfNnfa5Cb4l+FeV4BZ1sdx0nBejzNE
ThGmWrmBMsCfX+cggCiiNAaljCXs6mGDEN+dybBAxFVPDq7Xt910TYWwpguUNt0t7XUmNkDn/K/y
7nhlPuz3bh0h4wqlAXHUmDlHlNJsOCDYNwpMBASTW7KbewDIY6SSEl8DMF+NGlBzeDlu4fKHxFzO
gL0heGT4Xtb82oyEGWrgFt+fmLjgMjgtzKtjxlkugTYWS2PB+5rKtmfckDokkObMFOftSRt8uQe9
ucRY4tTJFwD9tVlnuwpqf+SsiQ9W3rXiSvWdcIwJDyhkHaqYVIW5SNBWIjzU1KUBHeXNu1hGTbnk
vjFQ247pquyNG0uG2eDnTpMUcvPyO432i225pJMh3eyuU/JP8brawF+FMdrSaGXRQNv97NyFWU7b
HVNpymvoT8Q+qRzpfkdHEWdOcrM9FL2YIVihgpuo4NC0cStzP4QhrOltAU9iYQR/5OBmqHG7HblO
W1q6DNpiumy4P+DVPBAH08bFkNO6A5DEBlpB8d5P2qzyPi1U7XJppnZt444IOB1MItGz0eWp1OUh
feppQDi+g0GuHHelXmb9RwpT87RyNT/Ys0QeLottn/stCFV4VGOK/PXWyHktljVY/0a3BZulf8bs
+FQ64zI521DKElFpCvqRWnJFoHMSHz+43sTr5sfqwK+9xVhnSl5A4y+mLeMMVtwoHPxx434V9rpD
w/PZ+OrlhomnVLKJXhhP/44KhooLRRyRlhDb35CJxcM2X4tdBTWkMCxKfswF1fW6CVwgSqLoEA6l
0J3WRnXN83LJiJd4UuN4+NKWBCQt0N5kO2T38U50WxG1MgxYkr+A7VwRU+pcBQlSdKCaW0oYkmlJ
ktdAbL4SAWLcxMxFt3waSaspiFZrpMYtBiNZYDxnATHfVXVwHHueMfDAPqx/NXOX+5nn4YqKkkLB
5wdLzJo7IkAhBT9C7v+Yjd1/jFvV4mjkQYeiLUVs8s9yjiTLnacuViG0K5XibpRCXiRKCnJLea0u
PoSFOVHSsIFYtrODElfYrSJWeFDGfXUpvP/JIeB0AaEsz+H8KKDbZUNe75ltjVmZA/F8tk7GypJg
0wLGsMd5ASr1knzyd/3kt+2StDYq+q5CE9hdm1RKHoJRk2t6n6Dbu9wSk8wgi4YIVzG5QKIrn6kJ
8p2pvPqrV9+Tgyk9AxgHLvASIT9qvzUjB/OPrX0FbutOEotzlWffmob3XzhtUk6/fWgICrfGXBvT
MtSoz+w31KO9BIUfuvKxZ4zH14+AgRr4U2ciW+q1JqIIKdhYAnbw+4zM6YnXxUZ27Cc1GtzgBnnD
mkVZISVJn1Mlc3Wlh+Hp4NN8ZsMDV/CG6iAP4ErOjgJrrhPSiJeS+VpVz/5X6zJpykdGfS+w4ZY6
1mMsgtx5fBgBKUSv3ZMYyLH1OG7KV4n/BdL3VwA6+3xLR2LCLFz1APJwh9ZDv9MhwgK7QBAWDOOi
PQu8YYghMDL5iJTN4dbktsHX1gtqS8CFBl9okpK+5Xi0B4hXv/UnbCs3WZ+6yB+yzIWQoU8boS/L
7j92Yo3hXMeUT25RUD37fY9HxGg58m/daN9/NosyTn0VgjDHS3O/2U9tEOtel2FowgJLz8XUtY6l
1hSaNn0wo6S6BUoZqYjBxG8fzlD3zVUhCX1Z3RcKbsQJDWM27FOU2PKK6vO0UzoMPeaGoBYCEDqk
x3io6mHc6hJw0LgGM7lDxurUEnSbyQ+WVMIQGqEToSq14gMOPy4rYiZn+ku9MQE0Q5nmPJbSlEhn
Yl7q8DJp2d7u0bGFnWdeLozm/KJ6cTjBJn3D5/Lfns6+zpFLz/NO3dUuTwVl04thGUHs5zRz4B1+
d82p79TcwuCIorugXOFtDVUBPAmkSh/QWdTIPwRam6mwt3/2OhTEzS/FhK02b19ra9PCdDHtm9Gc
KYxbI284X34wo0+5Z24b21o2D2ltFg0y/cQFweX0pUprjZBmPodnuq3klF3mDrBxb25jZHScnAGZ
oNULdHL4CTVneDslEsArGxWSUYEHzwTgjMl85t2/cVW8Fi2gy0ZyFvNolY0aUqbp5GaGFWVU2YBS
cQ3MTs6+RBX1mh5XhxPxlGktBGfilWwxi3i8Jzf9uYPkylKlP2Vl6ja9R5eCQfvDuLLKd2a+aNe3
CvGYDqyOEDDhz1mYOBzMl1wOylK3nJ0bXWQS4eOoYj6DgExqDNCrsk46O/7gWRdjHv2EEs+nj9Gg
0QBXHCGuelB5tRmm/VMWjiW96XsvG8uNVRb0dGeLMY8/k3NAYuneFshJdjktLIIvAja87pdwJTFC
cOA6/6s00mMtjUS5uQkcFRomZcYviHmokFzFPGPJYhw7C1pecDZnmHBQx7CzWkoz9ir6/97pmvnD
hmzaRxJVhO75F46ZWpNPSxkiC/ezl3d52g/2fvjm50vSzyIJ4vT5vmuwc8tJkRbYrYt/DnUsTYI/
BKFf9D5gWK1AEGBLjr4w0vehqn5HPjzPEwrZVx+fywicM9nhQS4DWEdwdAs+E48R9+5Vd5dFrmSe
MGBwnKhSbpt9p1wpXPnFctW1sE8uL2c1uZGXh0TQMp4cToB8atR77X3DGojH2cWAI12v0pDwEQGL
uBywfzIWIBkAEwAhzDtXUfohDWfpeR7HJae9yP7Qs+p9AOVMjWWK9UH/hhNIohod5DbC/47/Vszq
fPIEkynwN9Kz5I4Hoa6lMyCVjtuz0cEWq9gi2YUQ2VmyF1+1dELwkhg8+U8byxSrrZV9ACUKG7UN
EURKTWoDvf3qtei/56oKlDUL50xw2SPopImbFnT37Y6b5e33ZoS0emv1XGw7G3S2Ju45FZlUtM6i
oX968GqxvRz26KHrAGUzGmlG47mDC2AcQZ95nHl3Rex8X2Ly7KwttNe1bcKYyg1VSPRJuyn8cn5u
hxSVhfdcd6T11FtEZlMUgv8PRN3UHdbcHtHkag2oaJWjm/8aUjCqVdWGywhAfkGIFm4VwRq29LR7
8avn5eeVzFR3vUoz65HqEf0f300jCAAWY7E/8sE87oFdb0Vi9jDdbXIn0GzzfuGRMPYHpOr6Qn+g
6CaLnh0H8aClOIefgbIXc7/g5qMJoiJE6ZLkBS7qkFBya/magpy0Jn3qZc1XZE0h4y7JB/H5UtmL
6UidrSSa6m3Fu/7IG6fS22JQ8U0Z0wslADSDjuTpm5T9JJCxOoAqd0UiYpQqKp6acDRl0dLBqhgW
w/Hcau9bSmAW2hYkOMHnqPWWtZ+eWtiw6m9ZxWKZNaSz/m8+etn0UxtrPp0vblIqYtVGlix003IS
XkN8do9vmFVbeqrk8XJNvxcdocDkh/RjHKRxnyUx2PgnAQUkksPlnKcs+FGY+s8qtdlvWUOqBQoc
sTjRWqVb91RoyRMO0flYbAm+yPwkmsNN8QI9PiPIv/99ZRW2Uni1XlJvGWjKQvPq59RzzjZdpFob
AaNN+yD1issJhLeL3Bm2jI19/HOK7g67YHM487+qjV1CK954+UKUXYCdCPkAzrSiXe50VLsfiUpF
8yucMzSZ50Ci85hd/DvgXwioDsp4YTJvW9+52sv0RR6QYk3vDRVzvEPdCYE8zYSIi8ggQxw7v2Gu
m0B2d5lbUoG84887kLBXWP37M2OIqB5WRX1FPbx+RIz1WocPuDZXgPCk19vHHT9vzfjUQk1Eymb7
57om1yr6raJgG5+X6UgCIgCktJzAX92BxxjfI++RbVppFgNFZPuI+lt4m3ugL5EgKqXVdCdS4qf6
vGdl5OJ1EfeavLDOyBVHu/zDKRUBs8loOnEPtBD5mJ7L7/qY/bXfC/XXWVT5+noaMuwJDH0nfjfW
XEIRlIrAwykeuPpOwtv/E5VyG1wFuwa9qcLA+QW6WiFaaiNqqp9aYXGKw6BXD8ibMHrosOegquIW
XC0n2i53yELYey+I8UPNmY/FnmOcq0C1WNHg/koZSJZ/KKhmBLR3JcfGkJYf3Ddpgg5jCfWDdLnE
GLu55w+w62Xq4vKTY7PhgRGnfj8k1Tb6CijZSFXLfXTHzvp4jKgH4s+uC34bWQf1ai20WmyHTq+M
s9iJ6yl/4GVf3+1OtWtPOMwcJY7UZWnCFP6rSDDggKExMJGoBHjr75WslqBxFcVw/tLw8Z0ZtDR2
BPXV9DgRrfQK7X09zu56YdBDhm5voXsxz7gH63BWNs/ZyDnWnl6OkjY0kQEzXmrKt4vR0xUI2Pit
iGQOvcCftZ5s/SVbh1WSAhaYjkyuKAAnNW5OjPGEts8Tg5xD8vrBA8UksYifz5g9p+G1WXpG97kH
Hvi844Bo6CGgaLY/aup7RIhoQOwFZT0wyEhs+fpQu+hJ6aQ5etvJZlcarulDZKPjS1pisL+jhUaw
Y7UOZ3bhRTnGsvczDKwhgEEgoajIxJby1TAppiBbvwW0iuiIAgzNR+8Z5syjt7XEL3Q3j5HPR0oJ
1t7NO0EIzdPUTbXrJaEIq8+Bpbeee3YhJoidHMt6O4skyIvGPvZ6DTlAse9y/92Z+g068x3NT8Ry
hEF22lVFT11trY+4vUo/k5mRg9bbxJw4dm27GASlktkq0F5ziGsr3UiGq8n+XLeBXDK6jcQwA0iK
S+jWw7thzdwfzW9iTLRv/SR/LrnUrm/1xz7+DJIWBH0LxMs3YCOYemTFW4CgJN7p+VRAPmHVda8C
Z10dLddnnk8/HXPk6HAgHVv1mfk74VBqVV4/jZzqTROjTFyVOPDfnODH9WunW9ugn/BDWcgQh16c
37ACu7OP+pWBt3uSNR2zC4acQif5Zdk7siy8j/myubsrXlXjqYhSLrk65xb+ZRcuIpxbRykCOqdv
eATKx98EJvASrI25QP6BMKgU57ih1yNoNFq5aX4MPba6jiqeVxSYvJwsVkMSsFXccdohCnVF3KwC
QD1QusbEQO13e1mvWabIk81I1r6eLEhmyK/y9p/a0AvueTspULVqonQHA7AanSjAdRcQe66tLnU9
o8gW+x5VgsJ5CcitVTzkC6qGBCn45TAerKeK7kjOQjW/11KWWGLLw/Cc8u30fbb0Kth3+hmW88B2
FLaUl9nBXXjXath7V7CQNjZvfl48Um2Cyt0fhxjZmk9htrcuxtrqsA3OnspmFGnwnhuwgULd+SpH
IIl+wK6rGZKGM85wtbu4qD63Fj6fis8p+XsT1ZfdCWXW5IOvNQF+13ZKmdpLn85k5qaq0YF/VvuU
M1ZHpTMRDTCSJDPgRBKFAAQqRsfGfJq9SmI2mfy2hm+ZnI3+LJ9chkn5L04ARwffDQ+URrWpljPI
VfcaH90/3Zc71gKngQnK9DOkmxAlB9LwuhqfH3t08mS8Q7L/Osn1DrqFN2vDiVfod0XuaJY6yrMW
dD6KNKRo3eK8Ai9+vltum5HZsKimwTsm6psxBOhOmC9BvtTaeURzHuHCJv2okuoqLUws9gCejWIq
0QBBKLuYitNIk32TG1JbNixh13zukkpowE0Q+pltKt2QbiwcHI6ToAByBZYfiuyFICAgQWHnvWMH
e2hlVhjeTZa+nGy4picfcF8D+WI3sqNe6jtLH0Z3W4Ll72YxxMoWAEMQiM8Z3pIEd/4D5kEqJHO+
K1xh4ivH7dsxXryv9CV1trSVuUolo6i4P6rD7V8Z5gTDsA1zmjXDsaR1X5hcgdHPakap8YNQeg+p
xjX3yQvnms1JBLvmeeqK7/napI+msMgegQSyLkN46LOaz93MfD8YvPaT3cuCQI4qwjy6h8lJ3Vfm
Zic5ET/HOJD0kT86tpeaWpZYkKNQhPKwIlSPNpnCre1/aiVGtDel4Ea53jRDjM5AQmHamB8yyDUQ
RRHR0XlxRFjCRjsiHGPev3HprbWWQ+xEwvZ4yMbA8jMwufuvGddpG3LfQeRmO4KRNT2ntr15KUo7
gWGWPzrs/+yEpwcCale40DfjBk0JBXvPzja6C97QfdL4heAGxOfKckLlOpAS5StKtCvli3ANa4qj
eJeGHxly5srIFKkIvTUXbrN0qWV3IKXxS9VAcRJb85vI0mh/nSyslZHJ7DJzfPlV9iAzhdAUT8QA
cVkmkSSoqrYLjO5h/qOCWs6Qevr9siApW/jQwqdQ27gT6urVMcP4DfV1FWeLmoSN45niH4unkXxG
3QxC7+aGtu+7kXs73L3eeRfJFvEQTwz6qgg2XYxwNv9mhShf4YWIudWM6+odTS1lAeAhIVBmhqbP
CLpGHNSahRGs+IGxQOC96ktGyb5zDtbv9PEDbgdohqvsmX5HAtA8oZDi7uPzrTvi0QaNrS5dtNPN
yzQz3pEwcA850ioyttujm1xE7jgevY84xqtzF1tPYlUurJWJokQawh3yUN1jcRktNapDTlncgU0I
FsbNhB5DfTbuQWAX4RfRVSbHZlxJlOMgJEMK+SMH98iBVK7VYnSd9mkpPshmRjwzU4McFo+0LD54
UQQc9EfiuKnc4Wch3idWVLmo1ZlX6Xj2QJdr05VwDFQkC9kN7LQXC757jValH3wZ1GwM9hPo5L5q
mAz28UVQVzgWwKyhHWjcNrh0OjqLHVzZXXh1WeUFUkRmtVF0s0kfhK8ZzJI4vXyzHSVH1ziq21Ay
rZLwR+pmi14jYbU2TA1cG4QUpkycvqleQ7gJ6Ou76zdRD5soEXzPK1x79272Sa1BP+Wszik82yyu
DY69VjoxrySJhGPqxdKwDfdK7+cQ6J4u6fZ53JR+mQOTbSIh6LTBC9d0K2dAkDzmIfrNR8L3Ss00
Lbb+kGpHm1Dhn8+f4tnWyB5tIJvrbYAQw0kFHpGxAr0uCutbrZ398KZfqsawcJEPMO++O0G+p/LF
IcUpKTU3LCX1jgAyQpec5+xJ1eQWfpLy5sCg2X4Maey0IK4Hdo1ULx0FOUXwsFHRVUVtqnMdr8fu
+YesqNbgeGnxRz6GT31i4/LDVjSFZi/59R9BAJmnKadn/qxkAZcn5nQPe6jfkcLLi73zsCKVd3jA
RtLiHQj7Glz4C2vUbXQ6tbz4qVV0x44t3cptF7Yz/96csNLDhuwEBcMAdQiwH3yQ6soP2YdBzsn5
l4hJcQ2mXh5PAln/EREQYLGLUghJhyk915/SiJGQt/bns9k9qlFNWJatQJMlKNEJ7dOO7FgcQE/N
ncqHJDuVVTGKL8TtUGm4ZyMe5McuzMmQI81ei9IBgsCQ9OhbEPvU4KrqR7+NWBgbND0jkGvKSgJJ
S46RKolk1+ueOqSJ8PV3q7pgbbhngKZ7ui7oy59Xhd7rJj8thCBCB0zH66SnI8NXthkZ7Gtlahmn
Gc7rVLHUN4FKLS4Jd2A4X3mhquS0cMT8Jm7UGLLcGyq5L4cFh4nbZSJ9zz8sj2NssvzpxqITuhKF
rXUccHxQiYZ26lUXp2glACwquSGH3cTkIRKXDmMT+6fE04y7kSukTpwpeWEZ+6xbJMTeVfOafi0u
QV2oQfV3UFmfS1RInCFXZogIlotWwjKNQHYIZUNtspEkN9ryeq7IDHCIIj94WkbgXN0DecY4Z8BQ
6nT3d5cpnwDKJX00DWTPLU8m5+US+pE9aTCydbzjp7H/LWXdomqMC/ogiXt3qXx4NfmWbffFcaSr
jSQ2nuJQc4Uvt35dnyCUEFcVtQ8hmMzjU/NNNmgx8R4osJHYmAeXdW2cMjCbLD46tFZvZv6frwZb
KondNANvMe3rnoiFGa4dgSh9aGgIYkfqr6DO/+OC3byCxToLMyfSLsIl8Z2sXYC0ADMlILRpvRNy
+qaYCre6SYepviBUMZgWTuF0j6G10hiV3lN7weIzlPdJU0SYEuCOapzqlHsvyECiH2kiNHz3VOdH
grI5VJItlrVNCfMapmODOAReTes27sfCuNnGFCKGm1RR7tlAq1uu7WMBwoSf6+lxbWD4D5Ey2Dcf
0tUVe2mZMBHBKibQd86+X99hSWf795E7uXdgtG7YL04xPVG3GUlzML0WTySX7CiP7ImrQ96wfJdL
e7rDxNZhxJEUkhOMdCkhqrjNk5FYYV7lLke2mtiWY7XDqOQ9zUaI0UAvRhKd37ekYuvLSnYstzbJ
ArjLBOvdmne/3JlF/tHG5QsHhe02hUHjSTcejw0sB1EF8pfKNb1Z/gL92mhNx6Q4i/ZuV+DcHrOl
1laAAu5EuFy4IO43De4JQ88skhWdPsVgtnuZcZ2m0qRFUU1Gz/6ffZnT9I54xwE+XQm/IN04M8qs
AB/YozyExrht9GhEo4NCnH/kHknMn60V4acBPE6RXCXwlG75yml7N0A99AS/WRpw389WlTXF/oBl
5wvTm+oO3lgdxPPlr52t6OHkXb/OrPd1+dzndPMx4/nSYhwPAld74Mory77/sGwQiMM2AlEqOlQ2
qAB52A0GqRoeAHxjRnmQCXZPtBDoi3kuWc9uzDQh8tCflSLHuqVwV+7cLc7f0W+9b3ZZSosFvVfo
hMrOPW0CsQKxEUecDkwcSjJ4Fznapg2ldcB6UXL8c8fOpv37iNwEOaE/eBadlm7mygEWtB2qo0pm
w6WHx57woNAeIKn26NdyfWvCzWzM0GJANSDlxgVwUPiX82t3mxzhBETVnVUe9kpbm5fSCAXPSmEa
oL6hCX85Wa3OXtf8NJFJInMOWDJVgV6bTEobrQsDLm8RRKVu9P8qNld0Rt/LK0XJ+pdPAJ3htZmW
UAEtl1O93mL4ENBfIhKE24FHRVSC74tlw9N4zz2TIIGWGTzitlyw3tMBLfNw83z1qIkpkWK9QATB
ewHSL/XzRvdsX4OR0Km2sjlrXxqtaSw7EKQAQidgaXVf/EGVlvPObjRLjlb+HeuqXLIZeumf79gZ
xljnXVo+jNjnqduMu43C5Tx0XdiTHeYKNK7cbkPXA7Rn5B0dzlTD4LcgBS8lnIeRKFQyCYWbb6ak
wF2QNAEaw3IuI0E6YyGzWwyUYy/JzSO5Y944635aHpswUI4u/an7iT/MF9irA4Qux3FAzpJQC99t
lg8BEV4356tbOGuvavyk8hTVnIpBiFhe0rM1283jrVmhNwYuQUtgUo5qv5J5mHLlDTouNf0YOL40
MS9eu2lurxpjvP1oZZD7gX7uFJZh3wrN/q97+48j0NY5ocSYNVmUspR2UsLsLJ6p/+bhoVnadGYw
JmYdNquGfFRS5aPEKDnvmEQHU3OLOnnk7yjVZPeJ+QIKSqwcYcSdCtiLe+/WCGDdCbmZSKGkYBVS
oiDXgGoX/KIlVC2gRo+SIwbcFD2dJEFf1VIT/BRmvL/DZp4XiJPGhS1IwL0j/EYuwciGCSdp5hrv
Uo+PcQY4LSwq1zBMYsqXdcogy6M4NmD/LhWtGMe9rECNdSZHY5YkwjkN6Nw8AGRPh2oykKnDRalw
6+QVTUmePeu6lOMpf6CC3apJzNRiQWxDgj5Qe3uViS7hC3sk5o3BAJvLSWbZlk7345WKxFXQbCkH
pfK04pGLnr6JzwwE0JDSnuuvZSNCbAN35fbOhrIOExLEOe81XzTN+oh0op9mhPFf8PWfqBBgi7NS
Zo8M4/ZNWmSQRYBjUzFkuU7kHcrO1ZZSIBqxLxG8EXeM5JA0YILsKjKoRH9T9KqeNudj0KSvsxjb
AhFOOO0IZfG9VTmKNgMLWzFeHHqeaRZv6wNztAxstJuxI8dyOBzA2YG2MsiuTfbtScpKoeEJPMuq
MnR0lPoM8ZkGZbD9qQ8AMGrNOQi6Bq8cOuM3pNaAEchW7fBICylnkSnOTREdsbHCfusQFn6wm+Jy
dQtF2HnQt+zLPGnWHEZnrDgQWlhheiAOth6nnCsxBkxvO1PsZXP4bFcby5GvDsxuVbYgVr8ZW+lD
GBb7CWKRYg5JDoMiG3ahfuUA4Pt/y/v3+DXzYuNFFwzaRP6aH6jbFHcXPH8xzgEMj0acfDUOqrpF
c2vDr7VD89aAU/u1Mw1VUfqsO04oFXvin94HMWuqG/7p7Rw6OTpJyA7FMWksefqSsRMTFK0yeEEp
AaIv5FbJpOJKu6QLJx9E2BK+XnA0K3XagluJ/gErGWcqgnGEvEW+O/kLxHEws+DoXip25n4UCw44
lMIFbems1g2Vnx/DbJTN+xpRQOFwRGmmI/VsgKB3Oh3eMI7DSiio4Ftm6/arvrHe2xV/73FR6/31
okmxXRq8DNJU/WMhmN9AT52jcORhA9921e60qCp7vg73PiwFFiDOgsQHM4F4i4B44klr2rmIzK6J
WaVxaCRapGYM865/tWQjbcOW3K3Wfet+klzG51zwihBuj94tr6HhAU5kQRLiQcfuxNUXgmsELqaR
5JWuSLmihSolerDr7QrTodTVk1Q+OImiBuCxawNNOlgfwubmyBCfcBn2Dc5JGORGFgqbvBYgmGQ+
DRw34lMiQN168raij5b+hjTUbRw7ZyI2Mn8g0Dq2hDXAhwaRy9nbkWpapznoYGloz9zCANmOJQcb
Da6oSu54kVLXo+n4yMp8KICdm8NO3Qo4zUskgh2rfS7UBlzfLCDsLHitJRvGMsasW3khrTj6L/4H
OHtGGTN7eq0YMl/FMNLF5FUOTAvWp0wOElGgxPau4uTHaQ4zMXFcS/T+uRV2oF7Vt6P/AIGtWrmQ
ktBzROPub0b5Ak5b6ueYnJQmUL3yprsim4iXLQajVDoQHoqr7W6hINdfPuZmY8n1VNdNwdTFStuu
VnNAZsNwrVG58tY6DRWEYV7ctE1Ec3RErmkGjrAWQR3WsRuSkcmwsN8kdq3HPVq40sgwHKFcod1g
iUZZlqp+yjCHPfmDjxESZW0ehTLcU09OHQgLvBKhdIVA7CG66+eEMJCAF1fHsRJoAu+Kzas7Cd3s
2aMeaIgj7Kcp8QxS675MVRrJamcMzt2tcpAR+GT19gUDHAaPw2l7ahTr0wTMHHI2bJvd9FvoAwXo
1+h9fhfwepDhG1WHZA8MGQYJGddOCHDsMJcXiRvBd3ivj3MjXRLz8qDyC8LjPnTq8byvzkSSKWCe
+ysztZAcOO2GYCpNR8bhDjQqWG4K9x6vVpYhUDEmIWG+C5gs0QgYbnEt4OdxAhHn84a5lUQ0NOa5
Fby4SpQrqXKay4kYhCuk+aXAzT6BcMsDtApILNWoVTQrc8DJb+zThulN4AWB+tffC5MEmscLOho4
6Gvikqsj0YfYi2rcaE+H4S5AFi1/eRvXX4ZCr6hKDDkcBqkMqCe3D1BkhyIyUYWcFz2dcP3ynsZn
ULPmIoZeHAAldVHJksS+EKI9CdTa+I4fbs0cYzeWLcsVBHZHR7Jc5D8lzah/bN3Lqkc1gNhyDfGo
hku6LRaravinp17VAZbsGmujtzePUau0BlH0iEtWzXgoqa/gjnc8Bd2zrrI8KorJQ1GoMjalSP6V
+qeI4svbyTZNnnb/B6tLOo9Wq6M/2TEEDyBNmtiltts8qQajDZdDSrf4HHytsC5nOmA1muHxZGaf
4/Y2Ujiu79w3JkSXFzXFL8tz7FsY011lec3D9ieuKRcd1eN6EgLH20dsaRDfqZj0EeHbxW67RH/1
B4+YiDZQ+5Mp+RMwjjnSHiwO5ag+H/0LuEqvQ3vywT0wtz/Z9qtsx9QR/uS8KULO0/8Pb19Od5nY
ijzzCAz8kZDsooD+QAppj+AqK7VrADmAe79MB+Q2vMNbM0ojuC+GEgIzLKmf8EzGpi1TcMe5Iymu
YRtVF9dXQS3zigRtEReYmbiorf+NyR0+68vI5GZQQXJmsb+HlIvCeEHLzYxL++RDg4S/e7PGaKFF
2eqGldLKV2wlp+H9cbG+4btQ8y5uQzI4c5/UvwpC2hFFK5XLoAw8Yb2n3/nbuhsJ3cT3nrPPZuQh
FUKOm+lGBzkYXv3DcG2NC+6J/HOec4d1VEypx9p6yLlMq4VM549RtGMc7G3GzE+al5sxSeLh4hqn
+t2ZjD6AaszdTFIqX8IVMjaZpqRKSOfYvpjbx5ZkaYtVBisG0Zb1dObpiPgpnYLD7JOtK6rkhsLe
uiAbYng0sUWY+zJ1G1Apx0AcxYvti7TtReU0aMz7ZHgt4iMGjvYSRlbEMf4Iv9apENr/YRuODdtU
r7yh0WmS290VxGghiZ9BMI+PGFNt7pgBCNxCI41ZOTKdVtR1vwswfVW2LtvxJByI06XBFxbafjCc
7+8OjEEALwDyH+40/hlkdFaF0qumg5Z0GoMo7NdEsbcrNr4EWpLMwpse+doQ/7wYohuzPYXYj31L
0I2MnJ+KKMlxttl4/6/JVLnETtWGNU9LfA2yOOHPV58CW0nRuIgrccCwSY/+R3wJXYxrVOtQ/i8z
qVZDW2RjdOyEH26Ugtvtc99tFIpHmQ+jf1qwmcgXtQ/BNWepYXFYHONVbMTqgjYRA93+q6VeqwfK
hZksS/2/xu6FniZ16+Wu8U/vYRtUsa1g2E1BpZZYtMvW+e4zL5EyO0XBM23I4cZv1jsDkNpt6EAt
0983dNed1J4AdvxZZu2dpzYWdT5STYbpaU1ta7PdqloYtD8AyolNhw8SmjcP6xZDUTDjv65brYCX
gf3bEZLmU0QmvdTRAbq1xXn6Q2NrQyvgw8p+QJ8IzIM0g4LyyMngQ1wekKHtvnXuPSTwJ/wlg2d5
PwX1UI31WxRTtUjOj74DGSuPQWRIGU1j5ouoKEXm95iQp0YG0vIua8wQeFN6zYdlz8YI3D6kZHB5
FHQWFMENJ9aswtax0jcDM38IT8YOqoi7Jgt/+KPOm3f9FvAH7X3ePcENpmvmgUpHXtvdjSGjl8Vs
Z90rn97MzssthGM+j2Mu7tIQ2ayGboCdb5cSw+ZWZLKtGriM0OQHl5milM88JuejSlMMiKOjZdjN
xrFZ/4pxBuG5NBOIcmzuZ9j98fiCR459xrVfDmhVo6H/N/YjreVYOf4GwyI9vAID8JP5RlykspFu
uaWdNNw0l7JibXj/+a15qdik7xix57UtrLm0TUL/sOV+0keha+H1OSGRrBCv6DPwOXx4OKOt0RqQ
YUY3qIVBhfehSwYAZkt0rvaTAHehphve+NSbBQXz4o/gVQcm0MwZ1Wy///JqU1zz5X3DIEncdIaD
9alZO6P77viUjcrPQpIOr2KSHFLrrHPViATJMj+1KtXSFseyvy69sZlkByjFI/C6oM1Fl0VKpaXd
rWoA8p231IBvdVueJW1xe+0Ar2JUUmAERPgByaWdXuNT83wv3rHYg6I1FuHUJjwgGJXXeeDnkS6x
h9jpR7Z/AKzFRQ7YuXsYuOK8rlPdL+M+eAVce4Ew7RLt5xEwLwdrk7ypI8v3KibaFn8AlfsTR5WU
esAcvKg11whFEXm+PZLUw6lftkNc/gXakOWXKTRLfYOJ0newGoP3n5/Q7cDA8DWfuJfMC0Gl3MMr
OkBUH8LYDmVnnh2R3LlNrNgsUmL2MaZOt89zpboaQskctumbtt7+BmxSA2ZgDLnSDR8ZNoceG/O9
Y3BRlaTfKQvJYdczXxx94ik0IJlJ1DtaFkBU7U+Zyd7HFND9KZcelB2v7zqg4aeXyfsv38gHW42q
0RCxltT24Rn9PGJVd7iiOsQtLd4k7NTkiA1asHok5SMU1X5e+bhc0Ve7dLtkT1cMYPIHitezcL9B
YG9EhJZXwaSpOyJ2xsui8bysu0lf/g3f+JEQbFwVrjt+HujG4I5cJbmjnZ5gwKw9nWaZlyHCYeTL
0uqY1kqJQl5sFUd6a9OcVdcCs6bv2ao2zfmXyMfhR+w3HHetk5qClsWDXpg2u61I0ueZATv2/82t
dWg9/TW2STy39PEpYnLEx18OiCita9xxsoZ9ybaxf9bVfJLKxIkWUpIih17RVFihcCQqwSPs1Kia
Z5jy227m8RBuz9WXw1WX15GzC2Od5NfP5IyDzyFZD+hNqUnOAxPKDaF9AFoCtGDsvqQedGj3h0eH
g6rZdwkPjGBnuN1OY9TL7nafLKlXEck+iE5YaYARyedKiKqa9bI+wK/ahxSlyqEeZjvHpOpHhLgJ
d11xiRp9LXEJurrpXPEAO4CtlEox8GD+3ZeoecoTEFQsTAsm290NUHA8jcPVBdztyzjSSudh4LCu
a3ss30u0jxtmVW4rsXGTFsYm4Upd0TLuxwGS8FYER8vADZRtVzu/DJ57ZEVp2N8K62MbBg3Yzs59
++oGWc2pe5AxxDNrFOFX7u9HiE0gQYC8gW8KQeSWQxd5xxFqxlpx2e3JDK1utRjyV9P6w5hKNR6R
KBFe4ckwajJ54XTZo3Rh2HZ2+b7EhUW3b8guomzshP7z8gik32akS7VhXCgxhN1KFV1SiA1SHIEu
yPPcR1Z5EGfeHbWa6/HIwmRQl2cQXPZ8IlQGO/pov9aFV8RedA5a8AOzVROxhmQvaaXLg6Y/Jceg
QTWkhJ0Nop2+zNpK4i14/rcx3b9L8+hHAKmweRL4n21L35XqZiJpgZe1VDalUf8suHKVp5DjxGZd
bO0kEYfVW3lPG4pi7zWWeb2517PGVPlhMvH9X+QJ+IYrA65ZTzrZgxXAMUluctz0Uqp0eyjW74wu
zaduKbGD37bVuh+sf6g06Yy67eh3VZ0nnCzX6RHPXSwHP7GMcQJEh4gEk9uzSalWA6OfVCY0Fdn6
NsTwnt8yca/GJfsxWE2l0HdyDDWP7+m7uut4ckUOwngDzbQx3cDRzwdCWDV4jzGMQmsk6b//9kIT
VGw7naLqoeKb04yhTeVYFEI08iT+sTdYb2HJmZTqtA5qkbVKfWRdGtbi7vhPOdNSOH1RezXKHagp
SH8Xu9nHsXuDpZsPFd7hYguOtngNVgPqL27ZrWCZIHn83yA1u1iBMA+GMVPBF34yU7cK70XTN8YL
8fLQoROsW6IpqurmUjY46W67LsGrKI2Npf+uYPoAUFJquYpGZ9Iv+XlkqpB1WkUlk/i9ODx4HdRN
ENdkmIbewc2UDuMBhslXZNqMX9yKQJCysku1h5YH5O7ZUrYJxRAC+GvQSnyB+P82wFjj8vDY3BEj
1SK9DRaQnl7OV6YfXqn9xAXDhqfbabgIQjnltqmhXWQVLDuhmejBLPx6WuHQheQmpB3uj50HKLB6
UtjuLfqZMyyFn6BvkMqihZ8ZWefrBF+UPVpXQYASEsbNZryWQ5V3n6j3IxX8VaePXqkTLBqEWXIt
96aXnwQwBDJ5UBAAorNa0KeUo42nh7azVZ07LQYhVutNINA6ziMutQAWgUVFFKYf8wuzPSKQ70mR
Mcerqsau3mGwbTK4D26/sbOb8eVHMOXpnpI5j28IBCEo7B2Rxk4dhIU6sAPnXNJvPGccd05gfSHS
fAFGdg5473jKYbJpA9jhuPC7xy7y21PRafcg6sEumWvy2IZ8sEbuJo2W/9vZ6PXGe4fRlLdQJO2N
BGTofgyhNIDV3ETio4EyhOAJp/1QAc+xkaMPJa/Uhz8+zhdJ/qoyPJ+zvIssWAA1gsXHn42Q3cYe
4PgpNHTM7s6rb8OOzkZ63b1Fkyo6WVK1TrxsgT0ORiZbiB2blgyHGhkrkeAy9qkN5UTxmz1nlfrO
PZuWjQ5DnKPxXSOfmIz9xzIhi5RrmepseU1h32wHPQp4fFkxVoVpJrM3mKA9IHJ7OE4DZicFaxqR
TNQbwpdMlXRkrGfMISPrX2WNjSJf9BHwk6otOkjKIJvuLgg6ap9oy6xxbA3JIrlt1Ej/cMFCjIwV
OK3h/GFRBL1KyC83BzZQPCjfqeS3c+mDStclxrg71iDhEwyvYu2etL9xb9JKrspZT9b8lhUQbYXN
QwmaYfnbajp7kadgKVpvMjFAS3XU1i+hipIBg2DTPDLCJiMJuuNRRZPmJ/qVJE23XOesVEZg9o6/
oAsL+peA31WcY1Qhxc3PfhoL9XwDLt02LREvqvMiqZkTIR8SA/VWgkD3OPmHpSIPsteIAPN/2Cl6
z2dbS6k5l7PjIhDfHb3qoeRtBjotdArKWA/KrMs0FGszaR32X9GHKqYvn7gjWsuNTtMbTLRUo74Z
JQ6J1XCVLZI48tuUdaoEK9sed8TKKFy8POuhnBLOgZUqPuqEDH1RrBlJ5ZYiKPrazSFbJZwk2L4u
/rf8DXtgY36mV7GseZ0o/wBwKPgjg9kBo62jNZODiejmjFoVgxqFFBQE4vBIS6B8OBbgVI6ZzBBD
fl6d9kvz7JMBSrzio1vigKPfn7k4z3vYQGKz695hlEULr40sEQJYtN+deep8vWfALD+dXfeUvwCD
oo/zYceQFQkaum+Q4wh4qgoRicnfMZVlcY3Ed7sHugTzPrJrgwv1BqSVWxsqZb8Y91QF45Q7qrOv
YmYprqaJ771iU4y/1MGFoPRks9CLfM0XOg74fBwLXt5MSsTg2svXqKBFgEjwD+tZYpJaxH0ybjYw
YoXl5ACJQ6tscfZSYrP2x3Tdj9CiHHYFuo0OoDBD0cQrHSYVo4eLSBBQk84AXejjJ13U4eBxLkVt
2WPxBkoFs7mrUgx46e7qMtp7O3McgDPe6NSNecM/KVNgBbtHHKrwpjZ2szLmAiaEU59tkZVyFsxC
BF0XvrfIIx/cGeMUAZe2GSNvBKu0oSc3m05+J04XIty0Q5NYpv9G3usbmxG6VMMhayob2XZCa1ay
qMu0Pl8IoVnLV68+JipQW7UNdPTHURZA/8VSSRM0MaF0JV7V2efzT/aBQ/AShqylkFAHnPxccLMs
nnnjn/plR2i9CPX2DRSfHmdy540aZtLiRsMxmUVRHNPilbiFmefONLzRnweBATf+NIWBY5CmA9DF
fpODvpet/l/AyxrXydRaOLbUyQUma5MQo4W8AsFfdalJa6bkTsJFqED02A18Rv7KPec8YSzvW/MB
YFOqeZXpJEiNzreasqS4u19kW+Au0M0JwMsBm4YrBPQlDqB6W81832DWGqjfe/7wwO1wFQzK+B2F
f22fNRK3e+6/SvgLLCv5+yQHrZKcsJ0glCG5mrBDdtPriqfYQPmUlDpYIvcjmS+2et6fsRPl3Ls7
dqJ4ChgbEHaKE3h21c0tna33+7x/1qVS71+5SqodSusckiPNbVlZRclvrGQDTvpN4rkeQ8rJk4HA
bhE3MW+Sybe+5y2BCHTTLOPcYKLt1K4ZEFpNKyv5beuxfkZOZuMY9j0MVdAbfudyK8nbFCPs6XGg
79WxciAsHun3CECU16txiUWTPf/OxjIhmzHl3DhicT1mGHr83LWnfgZ4smf0YiCJxPfWTcPMsWD/
YwZEAUH7xUvl9sgdugD4gJrOH+1lqH46WQI3SeVYQCi83TW5fXCgLShh5IiIiO8EXS19M6tK8cPX
dnCyWZymuqB6+m7TTniF6C0uDdH23L3UrGcIZ1a0gUnsGVbnUK6qN6TJ9uI0AEa25s1jXnKRK1Qi
C0AQCLWzWhF2+nHIclMewXeygWx8NNLo06NqZMQSh+97ydAvPhxBL8+ZZIFQGsuvOstkTeAdKBoX
D2aG6l28drACluKcMrgSLDk/K1xJCFip03a4Qh8xPMPZjG6KAST0kJzwAFHLKqHakaVpopT93IOq
bwgHOmHqvfcl/0XAgZ7vQkmFv2SB1Mi2WobRP6CRVbtGeYj8018zEV3GiGs6Q0G3HN/ecRmaimm2
sGQoP8Mj5kiz+EE2L43+ui2H3fpALWLeXnmSdcWZR2Nkwooj0QZnSKhk3ujnLpb+0WCwebkmIaJi
VWbH4nR9gi39SbGWoSFlHZEigXsBig+EFK02yYU7qE+opnqAU/Er1pscHsrDbJ3y+hUt/I946SCY
WiOPeKySumTCaTTCsb0v67nyZZEkPpwuaaKTaqA1PRkt72OrjQCv078LeEQfTCRMNT+LfK69R7mo
wgO9/u4mmTU1vBrWcdPZxBjRUazZhxpsKTflh4zFjkqfFv/8nJbdNKXTphQIf11ZLyldssEnkh8R
6I0LXw3jLhUmCt1ioYZsdYZDjGIhu0muh/HWp7EZHqTjuaYreKYsXS380Z1JQFO9oEVpwk+gYH1x
+EcXqFoGT8lmqaKwhZKhMHqHqfcfjrnIlSFlgdlGPZ2ofjRzOGuUwX4sdJQ2Y4BusDmbk3pn7CfQ
2rs3t0u/OIggMWuwvhh4oroc4XLG70ndWu46TANnIPQ4yelebo41Xto8LvVjDVIA3nRclgBED+K/
gb8HABYzPo9rvsMRZKwZ6LF5sMx2akWnzTYkTQ3E8wIvqP7X4S5vHqKXEV93NJOqwEMCm5n/8O9k
EtRB6IJLdPSycdqmlD23ieMNVytZ+VXTa3JtxC++Mcis8YY5WgaekA3wl/t2Q5e2Q5GWODS1mKoi
cl5MO4UqQncBXl6//RtKV17djTSrKJKQ+YZ0jshVfZNZmZxRKqV5TLRSDQ1hVwyeQ+f12jbxLBbK
7IfsesPgermhkdFjJMCSV2jmJIZlHKuxDOFafdnD26Ti9+iYPRVeFA1xI1EoBI/XqKmqQD7BUlHb
R+IUEA8DR+Sc+uL3h/8S1eHUTFjf497YpoqUBcTAILEk2yLhBwG7WW1X4+e4o7XKY1qBRn3cuTeB
lSslrNaRXl5VRg8tgKjhHHvC8npljmVJoTAkO7IOTyyXBFaP8ZZC5Tg4M+gJA6SGOj3o/FVKVvkZ
+wa5twhnGOEqsP3cau9SHN0WCMfvc0uwfG85AA2MiwEWQJAsK4bxn94g+O4L5OOHtL27IKCA7jOF
e0QyoXhE0OK3N5yMzw7rZp3OgDmb9VQBFigfukI17ON7HO4bYkqkUIaYNnpEAbidNpIZJQ80JuOr
+1/NmOFliuM3LVEWM+VmEENJn1fQ6REWh5a8kFKOfW3ntk/Uy4ZMZwe++MaIxN/o4yv9DTwAY3vc
LAp2ZDB026D2H/CF8KKJaq3tnV4c30G2BO8NRaJ1yV9kNDk/D2tNnG8hZCBeVpoMwc9glJgTjuBS
6bqwI2gd4cOyRPeK/7TMO2jYHEVm2nAWbPVeSgHVvkKjS82e05KrXtztlVRCRS2cCM569E7kwCGX
z3CIIa2jS7bDPI9NYtW4dasVXAJWFVu+ZShM+C4kQjPqM5I01NudhfcyTpNguIHCRzALWYg3YagE
HJg7JbnFsNirs8+sq9x8zMY/ue3ntCJ37jXC1kuw4u0PG+BFbb1/LmmX0b7XnJLyNmVx+Dyyqi/B
5bjMfNu+TcfWJcv4CkMzdW+2DiA1BRTZJeFwPlgP/xEfno5gV6Nt86cHZoIli/sk2CrdIxFYMlqG
kZCkiDe2uHe+U6zEzDdErBn/OrthD+/ldGDM4rCy7vfpRVpappAzvbHlxcpFqQxDSfGCWhyah3du
9ihIZv+PSwlGEF1L2B4uzHCrmXC8PPUKUXBBZZP0/lHu0qGE45mlIKfHJl4icVzl3smsol2qrRTU
JpfwHAbMFNBANvk4pBmyk47UiHgmmA5X/CFzqzLwXNepJqLQ3Fm+nzBYg1yShZErsUffQQ/AEfbu
85vgNkhDecMD9kTslbgw5blMCDvXl0IMcmgRwYGLcFMrL0ImNK/3UwoJxrRbZ7bpBUkAZyJIatZa
dgqQmcTKYZJ0zzdz8B3Ngpxb7ZygWPjWPxTLTpq4BJDW6pR2Own4qRod8zkY5Sirjbp6PNxOw/9+
B3wzLl050KEQYwbx9XVg5Vj2g0eI+7wGol3fjcvph/igKKPaXDJUlY0Yuo8qP2nJCi6VWFfv7zaz
rplEhiqaqsIgot6JbuEwnzrRF+zqUBMPPP5iWh+Ev8CPME5XiRiEfXX27pCCHLnSoB8jzsmcX49h
0eXbodZagsQFxqigIqHmVkWV32NDguBUUwg9KZpiNV+rN5AMPa8u+Yp3eyLeUYqXyvnPVTWhvIQJ
82I/l2IvkfRw0DTm/kN3LmMymV30ou4sjAJ6+O9AyOQwKJqUVj+kUKDLUmsVxf9BPE5Qtjio0K2D
GYIYX0KHZgCKzYe3F3AVseLPuTZRA+yyA055lF4oYlWYSUyU2yPx3nWfcx98BmbrGibiqsjA5ry2
diJRVqLeog0Q+iEqyNDZ6pO0WDo6HlvRaJYLi6VFwYsQArluyyBLfDuD9mJodx5FA1z15thjPXZR
tkhDG88XChpt9ZMIEKdzXtAlxcAFVOD7rmNIgtzTExT1aNgJAfqZv+GcOLF+NcFCmlh1XrTG3kOW
k+md7Vo5CWmSs2BgiT4QN9pnkCDKJyDa5seCSbYsN24e14qIBZPWvzK8jy2evfG9RPJoBg/Vbwk1
mAKIw+tomzp84tpVnDcjfvP7fSZa8uhIAqVMQEMo8ttOKQyX4N0TtiqPTnm6D1biR3ASmkArNKEI
ZUDc/Irt63+Shv/SozSPamMbsg/ItoWcLBrxwPeeKf3xPxJo89DDHpTSqcUK8+8YlkU+nB9Mh1OX
fUccDx2J9gNsR7r3FWn5LsTtazJcBKfWnq31tsl3kiQImEjsXSGS5rE7Gfb/3I6RlZTEx0PWzQ+m
enHR2MsgBvBwX2yY4GeMzcA8t6UZ+KOn05mQi8QSBYDVs9CmO8xJKcEsk5jYJmV9QwYmslb/UDGP
wNR9SDAh4yunJQP2lEpcwlYxq6J2h4z8pE/CmmcH6rqYrXK5DrFrwhuO/bK1wgFI1d7TPUql85ut
LQch8u8OzLItXddVGVsP9CJo1mHDUxz6bc4HMtD/Ej66LjpNcB+cgJ7tYKzsQoanLI2McztBan5I
34/JTl7ePKt5T7XDeWwJTq/cO5QM1jLULIuDqk5XFckoZdWP4vq4M2tgOxJHhTLTyjYQG2rXAMlX
LZdTKIFDCgB6YAaa8M3qb/lfrd7vzLdZrA6WLqqVpmOcOsrTshNHtQ02iO4I2UAEHiXY9fnYOSOj
dLjyg9R4mkEmf7nDZBV7Io10M4u74T2gvH6DKT/V2Z3V7T8h3VUJMpl6v+vVnOY6u/tMtvpbfg9S
fx57JGgY9eaTfmNJePM/IYHaqM97q+SV08F4tLbs7tJSihGQqQNJmSU0CC/p7H7FDKPzLeSsup86
x//qIAfD/BP+cdbb1LgDWILpJW9j++TxPYzsBGySTkR4MZOE1TNE1Nq4rW0W1fpzQjpPbex6xImO
h4KlDUNiPV3LjW+YcmMUj/hV3yQ8rl2AlqmSc1yXlZ/xvhBM8iLb4ZGdOn3npTvbDbZweEmTjZ0q
nSIm0CJsgdEAIY/S4Gn3P7NG6F/+pgq6KAmK+K5jYvxDAFhVLYPowndXZww5ce1cGkmOEkiJ5CIx
2VFycofwesWJ2NQnUB+YDlkqVKk0b6LvpY+m32mP23ccOo3vijqecb+rtm8xUIaASWA4D3oYv+1b
ZGv/BOhTCXGljM2zazMwH2nhnjFfvGgMKB04JzMQydveQDCTza4h4ib+7ihY2ZxbPG3mI9N21L0k
hBQF5dMeEHMZ5c2K/X0YYR9neoWXrTNUnPX7ijcsD+WVAZEyZqtaH3eWsjngsAOGF0nKl7RAUUGR
Z/yUUN70QQNf3Kfaqhakwc6Qveapg10BaT9l5JG1e+lo0KHhUy65YHMk+E0TchbNQ3w1M3BWyc2B
xCQvyTwvlyMiHdWBF+JwE4rD255ie5oqGfp+b/IJ/W/3TI7ulfus2aqJOfaO9EuL7VjvqtT1+ENz
HayZzNOEvLiFsjUN1fxP4iJ7fgmA3je8ZkeDNac+jBglJgCx5/OdAsNg5gRTlch2zw9y/cjiMXz/
mcB4IfFBizy+E1ftMnegzFLXI3NwgqrJptmYkhrAflLD2gqnwaHmFJo2QR5G8Otnm/gF0el6dymP
IadShIjJKzgGEOozr3VzTo4sXRouriTZKDnSvgW6P80YGbZkCRj2OLiR28Jj1EcOhuTiN4daxx9Y
VOW9ZnA9v0sFuZ4g33/0IG7W/Yg2dlffhQTjhpVGwDxbNHGa5bTDziS2j78+x5LJXwPaRbVEVVpH
eNm5GjYrfQzOhWthIQw64WFvp8pVM9cE6iU5HVsZsTG9QFVMsUTMxAA5/FD/sMh8YSnp/jQ9a2f9
HtLRaS57ZXKbd3GocpAoZYmDp49S5WHQMxJ+QYDOrnyFjEwWVtCgdNgDqv9LrX3yWk+tobTy4FSt
4Sx5vCyc0xv2zq4XuLMOl9+GY1wodd74nkHvKaEyw6Dp2jBRhIufr++HXrKB4eG02DC+nWcbTbXV
utxVAssI7Vu1pzbMeA7KezZ5Znx+KkGkPilE+hBPPUkE/FxoIuxQEDZLAx2UYjT9waU3enzmglFb
/1guPrndygUcUrDiDp77fu2Imt3/JA7IG5vzgDfdUjjzlI20jE9Ku6sKz+UUa2yQiJucdnZwBAgs
NnzRIi43rhyJ70jzyxL0AESvO/qBRvsbP7rvSIGvhnP3SGJi+FFAa+0X0kcS1dxBBEI3tGd/HQln
hfay7nQGSiCYjlxRy8lqNcSz/4IoWQcEPxtl2o4mhHD4QhFAWUUm4+it2QtIkVxDw2Ikml6EeMrl
uPINrLvCnVr0cOsc/va+91XfexRX1pAHzAGubvwliJT6b2uUlSDOKkezSZnwzDBvmi8ypUtLOJzU
SADrQWtZB7LE+rkNb2qHCwcKxtOUzmWrMb0/daLNgsEqWLLTifBB1h4sLrFWsZesUpN3XZ2F946I
u72/at8SNn++SbOq7NDUIMTDLn04tM3g/gz2geF8yO6bhU/MOkyUYla8qCpLbzEPa7Teb8as6F1U
rcjNT3c5nbodz88eTaNhZBwbTNYKvUb21sYzOk/9l7zPf7XfNbVyVJOML//zp911LOkY2qb8Jmrv
F2chmwGpZbKkCmntPINputIq872mBquVovB8eabWhby0oUyUa5oVQc3JKeDIXPcfslTX5tRiytwH
HurQplcklz0w8s0ms+OPNnWfwZfWDT0f0/2Qmt9mMFJLkcDZ/ceagy9/YU+m0SDt73UcYXS7v3g7
k0DOEiBxNP/cV5vGW4wFSb0vsLFvtheftuvcNMbJc8JLsmDRyzr0SJtle+fNzudlzi/6EnxtUSN/
XRrGhpJ68FXAd+hsOh8jknaMgvbU+0sMCuknJhJ66csOt4v7sPtgBp0xf7p5v9D8h3dMC4N2nvM8
Jbz61DYLBRQ9fKWqA8MtLbwrGYMY3iwSJUm5uJUdQ+2aEoF7IjbBvd1XnX2w01/sQFaccaYpQ99n
CL1yLJB4j47Vbzjgy6WiQlHK9037kL6X+4mEtDuZtpMKgAJEp3CZjSDXBsmfBIRKSWUIs5wqX8u3
uinXSvh+pbFk0kOLt7OSX1P1n40jwK7xtdiszMqPE4lVYlP3MgSkeRhLy9wef6xIDE6Rf+y2/949
D0Uda5FLzniglTtsamBwUlSRSv/mMh59bN28MIu+UjGGZUItv5W5gwYrmNLOKrYrtmPZnik48bL+
EO8FmkdKirC7gTPaFsm8MwfhDUYXj1/GiORibIh0ZNXeXiVOM9KC3hQ0mTBF2i/eE6liUkL810Vc
NPMRyuWe0ayghwPi2obLPWoVR/dj79ussxpqdDAok6H1XiHWOHKqSCuZSeRycqWi4XgpsnTnr2Y1
rpGbUSUh3sRqoa4ScWim5tb+0G8GWDkTz+xhnWwIOeKgq/dHjMbTKjHKlkBSJuTPCL301rr+Oagz
Dnh9BsqLZOFGpn0B5QEEKzQ4Zas+y9DMwAJ1s4+ebR+EW9klGiwE8vTEsJrpog4KSwpSaBh1F1rx
eCJY1JQ0F+yduQK5ndz3hH8puJwwS2pxenDMs62JgPbqQ9Ils8IBK6p9y8CQQh7abCUJ8bYjm66L
Tjfv2D3IFFOipSaAVVqHwNwLXN6a8Q4lNR0Y7Kr8ZSoFl1MajakK5Tgui9QXFWHB5nmMsKvL0Tty
e8FqvIlfT64hrU4jWWSKqIbZhJj4X1Q8k4eo1FzoiRK34CxBwdYQ5216TpYQVkwk8bUZEh5CGsUG
ZaOYxqn3/hfljuvLgIULnUthYeP5obED8WGp58y6rxLck/aEP17cCnEp0UkNGvkmPspH77yhJX9B
SrWvNUg+c4n11R3nePyRbYpuR3beWRzZhUoLS5Mzt7f510ON6Cztyr5oKYmQS+5GvcokvbgLaPJd
IBK/+POjdCerqIkd7LlcRvydDDP8ThR+mUNxktwV1HbRWRqiICIuq6VdxN4MOBh7r+bKH7pKdtBO
pNSe8GsY1PNwp1zTZMCaFc4ikg1vqobOvp+cioVESwbU4ZCWAoXsGPVLMCdsn2WaEm4+eZ4nnKcH
aPOQzPYgQDGAkOitkw/UVrYzxldbvKaLjsc3OcXyaUa4ivE1frxTICq0l6ImHyDC2W8v6e65Acwd
9dMxhIEr7tpGpZLOk0NBKlVXcvT7MwgJDoc8ZOdSLnbBmhBeUn1jRZ6RU40k/LxOO+eLXU/Yv/F6
aNe7rI7yWEyWiIIx45onrjQvKUxLrTVBvpxui272jLzn0BfQqPH8TTJPKfXpCMaAw/Nn8PBRt2z0
JRug5FVJxbbZfFtgUSgUnHrna87v7wMsiy9Fxi3otH+SI7LL6sg4FM1jGsWYTSwk/PhhEXPJg+8j
1Eki4ji5m3MVMlnhE9CWOJTgF1pLf63KeRYU8UeFBj3b3UXZ164d3ZrvhJZw/yvClMjb2ORN1ZZR
ulQht+b0tSo9DilzKxYfdKrgs7FRa1iLPOekpSUvVywnE/8qxDIdewpaNlXYJnBjcoN3JB+AT5uT
Y3CZHTKpm6qF2zfr4vmXZSNzKSRIqkh1SQS5V6F0QqVcI1TNz3oYrhFTWvsBG0Qf8r9FysF+frWD
nchmBdreBjCWs5Q/ULs2sBaIyYN4DnhLa3+5l7lSdK9iQC3kVSgbaL1C1uYB/AFLdZPgWV6ct80r
aytf3au/h8lkWQHmPCSUSOLF3aZmNpw/GDnt7EPvL2/6SkG+kNyKOOrTtcXZmxAJnbu8BK5Zb7jb
POYwKvD4prl96Un9A0Xy1FrnNK+GIPQGaNtpnmEsphD1gaRtr7XS9uQch9UJZB3zAd4pBkHlJHO9
1Qg5Q8bszvGoOvjz4VlupwZAt2VES7+sKAfuNwp6OVeb0Feg4wQPzinIP10AQ2uShD/5peSnvyrr
AHYn+SaYn+b5wRqrCfm1H3gKHr0LSlCEoMa0EB7U7pid+NmOriJpRr4qJjtrQUOVpMJ61nsZ//jj
qcW3wpxi/ezU3EAeKjTpiX1CLAkzUr4AHy+W7kyH7ZaKdx5aUR+X/j/0zLfe4NbJwomI+QOHf5NJ
tZnF3hl1MZrUEO6PeKZdiin4b3Lvf6zg8K4YJLjC+A2x+XzplCzZuTRJ8EYaK7VLHLaZTjNPePtx
LApSTtLewXZhp/NPAofrs53EfnvZUQTTYRayVe9WzJi5Dj7n/8I+RPQzMlNm2x4SepAI9fP2Tzqw
z/u8eyyjD757v2Ck4pAcSEu8q2ptE4qO9P1pMqEy7ywvD6ujVdzvrli7PrfXPIPztMnPhPmd8K/I
L1H3fK4xpU6GzEo20xT26wWG/FkcBUDIrDVKv3Jx0EsiauLKN0t+5MA2XQ8MagsDjPq5rcKh45SS
5fCvVTLUBJCJVe2SPvY19tziDBN3QUemBmuYl+UgI0/3sQv6Ac+mvfqY5ChdGfr+HJRah1+Nt4lG
yDeHlRlyHyjbZnv4dIzc0V9bLJP1JsOLcgoM4Arhed7jI9avYue4n9oZC4SxDcOA2Hf/b3KvwiNN
eGju7dUdShJKW6f2mPIl15Gz/DAMLTA0YH5QyTB/ViyK06TiAy43y793SfTt1eM4oDgpnM11J6FA
NhhiZqZT10sJtaPhfZFZ2OXXTCUz0UTtE9UsHkDKAOYpxeD/CKc7S7bOGF7aHUN+c5kfNr3SGYjm
HpRynsuOVNPZkVntJ3cxrm6UIRLOI5BSVjGNVC1noV34DDKzcYOEUwlTOSqZXHcrd08hlGRTzhJH
HTSOW94RsxkK9Bd1vBGliMgvXIk+ydAzjweHLbeLnW6ZrnTmtH3xMzwGr6YOgoeC+FloY6KAyehW
hM4v4WST8rfc8Jq5FPA0dI02V8xx+vEZZflT4ygfU0z62KkP/khjoDNq/pawbyZLrOGobLNckzs8
Mt4It2Xm3FlsQWvwQZP4m8/CEtVdGmWUBykvsdong9mGL4fLrzx/eudD5hdR9jEm/Lr8AOwOQMEp
494liDhwzKpEnPIvovWQXsBOPFmbrH/oBDW//4nosbt1d38CWixbobWkHUEsQxCdFBUitM6sbB/7
2vRwnTr+QwhV3RuTL23Iu/6TbAT741WXKBJYxnl/zd1UFJeCoVWav69cjq1Ea4gQ7WZkDPr4I72Z
jEA3zAuaBptTOZhYJR4lefAyyLZlZaJZdpHR1tibNIS+7QiFsj+DWlSZI3gxrBGCQqB8N3DeVlYQ
TsYwFJ7hULeWokIMgkaSdDI8ssmtLHwYDvO/xVUMX8Uzg8cBf9ugvCYPp4bsS7QGCWeMHu1z8xaM
P0jeAaLBfsPPJ6mAnxbjzMFWC/G+uD9+gUKvqdgjNpeuRifxMsboZNG01ATIg6et0pRlw3nW/XEe
jHEaDGq9kdaxOH8PaoOAJFQLgARJVg9vMoJBMf5HjbQe47xTA/Uek7mWm00fbA3mSPqOkKA7GRPE
tp8zOhU6PXNHLwsOlXEeRiXjT2cMCe3zMGpjAXQ5kiMtKBH5yuNfVKrP1GH2ZaC4ntJ2QWEpTG5t
bhc8wwcjMtZu+KWVWR3TwklaEzSopVaMYXvSU0F+aHWPQRIfOoBPSxnzmVATNsQLDwh9SHl4zQlr
v+BbqKLS88dqI/6QLewnxrF5YNXjHN+wtGfn51vd6GRxlFE6gHzl9I1tIE7CwGfjV2+uMgz5dO/P
+ElMrM89Eh+b0KsHzK/dPf0dRqCDFOwYJXfwtwpNKhCZhJMH6AttdiKqV4gIKwCtOpMLdxVKuc21
l1G4+9Ql/fQK31SIfp1Gu+0yFWzSMMk39CWuDIFTCVD9NItmyuiK1bBuie9j12i6F6H03ojmywf/
hssbtfs3YS8OBT5eruN/mktD5SXdvreIgT28bmQu4OUtwO32YA30oGs7zoh/pwOBMzWt/tuUGxyw
Yd9ziSi3XMQDHSJZ9LJg+kMJPAqPk4YPb8AnrHYqjllqELEnuTfe87Thw2KnqgVl13+eFaTSIK4U
oFh9wEIcHOsNLn1zdoneyNIzK3gJ9QXF55/1770Z4d6rrHJLIQ7vYqQcHpqCmOmK0qLEuokM7XLE
bRY5tdp0z5AYnV7QS50VpeiZrO38q2EO+lW1+eRoOU0BcgAOAahTbnoLHhqpgcy3DpRyWb2cjmbR
FDkpmJcdMHMgeKn9QGgzQi/jX5+z3fFdA3BlomB81yrsM2TA6KwevhtelEstuE5LjNqsqIDKJzta
/Lx7aeSnx5941stIEjErBIfV+zSCCWwkpwXfLnuRT8Y4B+e0JH93i+tkukqpCs6llIHKV1hBNFK8
Ad00pEgX2yDbWiNynlYIciUko79CUauOx1Xkw0ZC32ca1F2qPlukN7mF0+SYciUbb2m31KURj0ua
OrCVyvwdShX5vJH+20xp8E5sATYZTmlOh73dzaGoodc8+Iq8L4Ow8gl+aGJgT7TJZI9mWGXvp4rk
2tEZrLiyZgZBeP86HW5XyHXShAW+DgM5EHzJZwiBpnfs7HAP6ROZyfNCFfzILqpecT2ST89vaCPR
uXIRIsz3yzQU1/c2Bp9mu+Vzq40UZSQc15lvIYBSwHJIRbYDOYUGLRdiLI/yVJ8uhElJ+iYhzLwN
XezfpcJ9qe/zvQPsH/QC6yWGo+jv1pQ4cq+HWkqCwKpNGv11mpBYDTLKIIPcrK+KR8ZZX5w682ns
yiW+tlSH1jTZH2j9kCK6MecWXmVBQGrpcrjEy0ORf7UEysI8Amatgj8uWrZpesaeMzjp8Y6kCvht
jrFBrwv8iWoLVv0Bpn3kxF29rYHWq5BjOjlhxnuj/3poF/tvGkaqPfRY5uHtpoXjq58Lq+YJp8uA
EaMVMPWQQNBqUiT8BQOTzobtpHbi1N9k/PPt99Aw9N59kI58WzK70d3E07TxjbLjpKuFixZnMzDD
c0eEbRsvqF8fyn5ex0E+LBUlUO0xSACkf3wh3Gm0myq+1V4HFKBosYPWbykQHOrMwnavgoglyiBx
gQvnVQaCOm82YErjTlRLFd0eS6QiY+lazZJ72+09SVE6MfxEJpqehweU7+6jQVU3DP+HwCWcou/y
WVaaqSyYSrF2Ls4OhG1pOG4aNZvgMcl4bgtD4vxYJe2NYPe7RndKaJJBszyGmD1bR3AJthUTdz8d
ttjE9+2gJYdH6wE5vmPGvK24C1ucXWwitEW/+6N5CJdDRPe4c1/4FTwxbsZ40dFWmmjGN/rxMyK3
Bh90JxQpXP7HV0Mgp1JPw8rc08c4Bqm21pSGZL/BwPo55eh5jRxUFz4VCayHfA7Uwuqi/yFUoRoB
cxMRhU+gkUymYISaL1Op6gnYFIlUYQKWpbRFX/HaWW9JohPCU7TzKzEbuuJ4in+MfR+MKXNwjTz5
vA3TtxGtfEtFuppPiIxB7jKt3DpsES6u4MRp2t8CxMEhrb5CkKYL3UgA3n1gwbCyxgpnB6gPS0/B
4BwaueYmcVoEOTdkJaw8L4YUfKnIrxVCx6fZZFr+KChJRLork9GAXNrHJPfBCpkrSS23Ydt0wFIn
/rJsOl7MVIW2Yn1HOOIm6K7jP+NsJ9VpgnVkPr6Bqoj5SOetTjoSENHb24ATbXBwWeuvCm7NbaWu
BmgyPhJ/vhN0+5oyDRuXqp/AW/7gp6nTWIXWtKlL8A+Vkc+WmkOEYVQ0YQw0WJ57SrMlyzGWElJL
BZE3pw1uVWZTi2S1IS6UVreaWlAabdF5TnIPNJNH/3hI9URYGde6ZgVKlZiS33BCHZdO5Dj2U6cQ
J8DSaXeVm1NHkdAjQRpW/Nj3/IbHLNE7wEltmEaQrpSiOKFT+OYYwbSF/GlJ2KZCzKPgv2SDDHCY
gZd2JCr8Cdbrrx9HACI60KT1OV+MK4niKpxl0XnsWS/Z9NKTlc8IsYJRJ5+vjzvhijsSpEaSmKx3
D849eGO757x3V1AfkGegslBrvwBxPFlIBZJmzZxxS60LczkTtlXLgtbpFUQbSatC1fVKoX9sB2MX
GboFChiuRVPczJ8d6v8lhf8cNuIOE4TD72VTFUClvr74WIz/iw7iZFX5n4FX02lQdhDIq4tQgEIo
nsEiHSh3avwobpbKfYsRQlqByQVjkMY6ZUjgLxvDrekA2rruk/ZkceXoiQxsiqxnLXZv5RE/98zA
PyV7O6WFree4AriOHtM7yXVAq+ddWLyPrT3qqlxyJTYGlFbr9D8Wpk45N/hmgX9ZPmQDuTYBI2ci
zf9wNHX8oJ0MLd+DtcFtlDz9sULc/oD/Wo9vs+QDmeufbMPTKKU6Dm3PM0z7aI+UOIkWRAUjm9x3
LUtpx8uuGvThVZ1/O4KUdQNL+CG2mMywoqW6TfdcIjr0TH5iPx5aaTBiYVbmlLuR3W8g2rBO4xFk
QU5a9QFpQBEE5m6IeppqpJFejNYWwcewYd/A+rIKJODkVItGjrOdTOQZ7oGb8RieFT3/bpv25p2p
c5D7+0x9CSZHv8C3KtEIPl/70P07l0m/n7Nn50is/ULtfXjXUiGCrSXYYbYqRQvCK9mmbfafOw25
916K149WTdN5eeCcdI3DhFO0Ek1+wnWp8+pdUAFyOrbmHqW4zebnFWY6sACDIwvQ5ETDRF5bpdkD
g6XbwzmDIdkm47Fz2Qt81II/XePFDefuw4P9fyOBKUsy3bYno7qIjCM+B02q98N8N2JfJqfD2RaD
q5yRGinclN91E2sIMXHgsNK2S1q6P8j6sD72HGjQz7vHm2HVIpUMuZH8SPrM0hV2GTMhYV1tkanT
7bPhb57U0x02gC5KGsPkq90NJ4ZFblLJ5oFG6NmXTJfuxsENpePgRXalcJJQ6208uyuWyPMGxwpP
4h9ZwTrb1Z3OAE40x6Z5r3gkfzJCTDhk9N7qcNNyEcmD493Bmkza/rLr7P0dQ5U9fHEFAOnjfd/h
yYXEpJyvGdZxI/lquc1yJ8rnvrc3M603WrGMFRAvQJokC4vsRGKmxR3dc/M4r7VhfspCvLYSd7BS
fpiDiUs/vYb3rC+LOlKIk5UC8oyaXFJCvL7v9EfYv17eJi+jLeHQrqEKlu1TmBZP8XhOGX8JQK3b
EDcaywPsh4Ce6qHb8R4aYBq9vya0JUtnAH+4vbHJGbfY9VSisdIiYhajJuEw3OI6gGrR1lmZrPFs
eP9xi4Wn7sz+/XumhV92ikLexNuvng2YngfIs1t7wbqQMUl0F+SM0ayKY90QsDekPZ0EFU9aa1Ib
879kJoCiQWK7yH9Fn3hUOE5TdlHce2l94Az/5AWG2ZjOWlIQUTbT7M+fJbu3OYgGWWVajCI0ESNT
aQQHnXOpQ1z5UhHm7ohfui6yjeN5FtU/O7trFA6T5+5XuGUA7Q6+MkU+ik9AgxgsKknU6VQ6TqXU
QOM3AFTphPuIJdLcITQh4FnWKqMMU61iBcUi1q3IZAzYGNRaWc8tFtHTkxRQFT89KhpSWrF5Op82
eyCU3IY0ZHAfAU/e8V6wWpnVamZRJNZBR+Wz7aorWpZOmbVoMJdpkHTIJp0yk2aGHnI17atapLTF
Bda0hQ+qPz+qibCrbampJ1fVnYnTll+2Qb4C8czCpruGl2d97+C5JGRDBmTkUndiSKxkp8Wmk0qM
fcmn8N0xp3BBg7cPclejZTtC0/dvZ10f+M0LofVaogEn6GkXFx7F6aEArLYETeW18Fnv7AEBhxr4
dxM45yzMIX2kQwwR9OwgBHEzyZpUw9mXDw+UBxjynButRYt8opY9j0BTdWINy+dVy5SR8Ly2M8PY
nSoghi/HKnq/4a6hYAX+fcFnAZ07EiPR9l/obhuikSkXiJhC+R/9Ww4Cdpy4ARV0IAkMs2v5zmfE
6d8NmAIg7UFZl4DuLrQU5t73gGbwz+Kom0jCqDeVJ7Bjcx1973eOflK0+8qNmDn7Ls4HAhD4DxLm
Ytfuh5q8jE7tk3IyGNZkyP1ZVIiG1oKUX8uOnhuQOLeLEAgsd00dXTdmwy7UrOzjbcmWpx6HyzM2
SoeGLm4tHA3UFn2Ir/JoMfEoUKL+hDiXak/SJGFsEfVoIt4mrbINurkhPWT4jvMpOyvTjIxOfBCu
aER4s8Fd/cfTSZjGYC88I6rS/e/QloFz9OiJ6rEAF3J4ij1YdBjJT8Sml+Nx8z6yqQkKnFXax1B+
gho0GOkhyB7o1qkynxN57KEFuIWqSxDUZyyo7UxKnFQ+9Mmd5afAwpxhOpFg1DV1b//3AUfo2flh
M+CrIlVzmTqdEZgeLzwpV2qiOPb7jndm+B5E5NE5NmHybZ6ku4sYzeCWwuuRT0Q3TExN9zU2tC/7
ZuQfdEVXpvlp8LASP3A5wQxW26fWFHuiQKxlhCASrqLQ8KFW6+UrNrAbnqlLCZ9gAppL8TTtZwD/
KL/j7gPvNFn2zHQtVAwfzp81DU/ivZEE4HeBjxs9Ofz0/uP1nXslRKGgzbrv8XkBAeqYX3CIDt1M
4ANTR1AsHVXUPOyGIAIJVkzvL9FsJyH/lrP0NPfgYL6PZKWsQLUYa1g1w1JaMFqrQ6O9hYg11OZq
IHCfw+PmR5jrDzvoDIxY3qzcoMC6YfqM3goeeVdfpcegbVSvndK8y2EKxEpf3UN7YkrTZVWMPxsV
chZvhBIRDxnPn9vs/5r49YNl2PTtTF8qc//g/dvb4smj2n+3UhHOZyGhEAw5yFm1kBMgCQVVK+Wv
/+jZbMWUcWTJwZeqeoW++mZfPt+lOwTH2joKLW3Y/oEi/XKytVbN6Deqatscq+AHy0hbLe3oUMig
wbDFKc+8BprR410twp2lKjHbMfJdDnBCPHnxtYSPYelHcThmPOLceLljwRmZ8m+4PhvoOlJY/mwi
s1Fy5cfpBbaY8Sng/ONuR7rc/G5CiaYW/Ci1HcTTIpvQqlXy+E+lixmkMJFE6gsUMCc4ijNpijIh
3fjeJBp1sUo4VvOdG2Qv13k0RY5fb3USG3gMLFLW2B5O+4zTs0fyEkTy6IXl16c9BMLiF9GoT9Fc
lMC9+1HpIJocFraK2+5DROciQ9FW81d8q94aIsXc+erNTX2/GK+X79ryQ1ocnPTd/HBqVSmfl03c
/R0x6k1a+5iUv6Gr/I9omnTct4aR9S2VOrnYNppOiqp3cQhJc4KGHHyqat7WvHJf4DvoxJS5E0Wg
2wI9ufOb7Wv2l0vO/GKUd1UIjVDWB18JsAF7BCXkaN9w+0JT7/YN+PzWrt6HG3WKbZJ0PZFGKJeO
YiB2+aCsaqGjjrFf35TiTpSB2qplcEAmens19eWSM2ocqDcjjLjenXVLKPoMBfXTpaZyvCaRr/OJ
DaXVl5hDGwLpnYNJtt9CVZHatrXmyLhEdGDcy3kL4ZUVFamMSstUWC2+IeYDt9O+U3Rp+kaZcmxO
jSmdnfXVEbDxg/7ArCA0uPdPCATh0hg0RU9twNWCTqi2ZNBnXdX/v3OU0PmaW+tK0vdhOdI8Jdp/
6F+v0BEfvGXmxZ5oywGFsReaQ9gQnTwEB5oE1SiUVkDIuX+sV54xI4BMNeXR7/tHnrcyFPMExPaZ
Lk+NzxiUNP5r14muB762p5utM1wrhQ+ahr/oq7HoxnW3h8+HsOMX19AvkznayuLyiC69UCzzyCNh
uR8KFfrnzfzkNMNwZAQyj7hvmvdz/sgDfU2Hzqt22YjZLaPHd0UaA/K4qyaGMz4Lj6SyqawMTOuk
o2ERu+9yiiBzsfAKQ7WqtKCRSP4MLVQbiOhA3enye68CCDqIlm7HTUHG4c7VpsqJuNGQ/sZqYYsP
YSBTX5uWvfnO40wcHhDG2O/TBBAIZu8ZEe9zFh1GRDERjIgO+HxHF++So2o8Zy6ZaX1Bo9T9kQS8
Cgz5llIrgvECvI47QOYk2BzF4SUTdMDEQZhnTTrP8iT25lGJf4PSAuJnJSnOTiAUvm8ZrQC8A8IA
OiD1xzr+Kl3Ext/AKS3qjFa+qn6oDBMFRQhPRrBxj1b7Se5b76zNpBcEYtSiPsVCOglVyIA3/xGl
2W/mJ4ikbJ0NOv16Jdsyz2/K62O6bKbi/woWJBn+ndD6t0Gz3d9+PH7xrfVztMr0V9pVw1YPLvwX
bD6NK1UcsTpPlpYK8OAkXyMqtziCuS2qUeKXvhWi/Kq66+nbMqvxKy+d/09DyPgU7VDyGHce5mz9
8FwqjDCVBYovMRwr3ajcLy1fciqW1GJug5pf4MDqi7jC/CYizhEfXfBj+d8MGPNJHZ/AYHJ9Zawu
7uLd1uSUVTM25PQpSCpi8gbncDc2kJQPo5r0dcGKdoogXQ/xviwWHicQ25vYpo9WXYYtHAV9j+Dp
8mHPUXENVAvyVY8vXPzju++ZdCDmYsPe+VwL+cn6/4jE3R7pFot2nH/h9vfyFuQJYYV9bithhbBS
DdWMdNZtF2EH4WaLAGRl+ouoUYyB7cf37WLi/1LqtnGpjgRbPW3YcIQa9CHBL9CMHw14Mip1C6Fm
BKtH4xcIIB+LPl4CqLTrK9DoHvdE5q+s8yJx4vQLVQUq6raWCwrxWRszpI346ZwtH2T7gQB1B/5M
xq4dNXdaPMj5t4PlHRvfcc41iJOQglkNkgatpCBaxoicrcJT1Rymjkjj2AplWTUKJNeJPEVX4MPP
zw2/ddOFvsMcEday2vC/O6H1/0M1PWMlOhP3oDVPza4joMYo5Qd+jcyf5S0sisest0fXvjlzpzTK
vLTn8i9nAPJ7jxfRhe7X0rXDpANmFhLWVxm3RHASF2o8GKtMr5vm8evUovp2nfv9WA9gtNnpx8KI
TKTwaBir2+d7g40h78TS0a3Cn95qlKoLpuF+lsOn/BuZvIdbEK25uyCBOBnvqg6jZqzH/5nC8tCj
ZvxnCPNxq2h5cJ+lRl5ZgF3Jt3ZtOKnQkeD8FF/ZmYLIhBkE3dy4UKjL1J7zgt3r4isgTlZscWcr
0nDLOn6X0a/XpixIktcpZ7gViC64n3bc06zVFD8S7mbpMorHgcbkyhGvWClTBZtJecfcA5EAAaoC
pI0/vZlorCBbS/bJlrMO7qglmjf9YGXZqMcOoEoOBZn9zm9MTngPFKXkkxxsPLb8G9wmRosDWsfI
IL+d9DaRT70D0MFq6MnIs5dvDVRZOxmAh+wocMQomu9TG6ZRVIIPE/5n40R2Luf4Opb/I65l4Blb
lvA55DMzQ6yug/+9hwzIk/HISNtvoe9ggf3b+HZ2OS1wX9HVSm2Fk4TsbsuU6JiXJ5Z5yHJZvLp7
o6omGMO1qeNfNY7eFX7+HTOGGf5z6NNqngbUaxxRFj/ZJeVjyvCdO9s5zCr5oxRUoQ5wIEVUUaES
HlXyVm1oCK6NNXuE4zDgLwvWPVKplu/rjAfLYlhzThHHYzDC6mtiIGitUPxhpHZ9coS8nqu7smLb
1LOnmbQf+KhyKPagilMVKytWg6fTFdlxpapuJxoo7ibVEeM3RRpPpSNT95g7wN9uIiPnBCykBaVq
hvohwTHmh1xhmr3/h3Ngsb/7mNHh7o4U+EJCMwOELUmHOwuMpNXAmlmZpuZnl0HuUAqU3P4wykmz
zoH2oTQJv72gZNmwRudABuXU2Msxccwdy7lDkV7I3edeCKp2dF3+N3u6YTDwxbQMRv1xd0Zd+0k2
/emM61DT6niiOguh7DKIRWl0nkiiuRHpGNueej8uFdFg2xcpoFX+PybPoKov1mHJNjtY/BJjPdF0
MkWTPumMYz8Ry4Qdi1KfB8JQ9+mkiSt1gGhUph2nBZmIrG7Stnk8+cGCam3ntaAMYC5szfLMZetC
GIprSxTrqM57v1wUisiPqgjj0atLYknaQGhkzs75WY0vIyx3B+cHrw2LweKZxpooV5MhSz5RsFb0
aWa5VYdskb92vIHoFTT35rXYBU0eTbdGfCgfSrq5799l2cVj1d98S4cKZrtpoWZtLVwFQCY2XViD
AjJIkZQ+NjlJPVM0byKE/uwGcfoSzLDuwCcEEt3C/WWPAKzETIs0Di8T+OSOxT2fbcWgb2yEFt98
MKyELl4/fl1La1n6zd4IsqQXuA2QBIgznDfg/qaib3eamC7JYp0j83C+8ejLS//kBpPmSttg3k2x
7jtkvt23CKVMUQNYFA67LJkqst++fNDcazRWL+ujCGSkkhRdAMYmDyHhvSIxjff9traYTuFvDYoZ
pVyOh5rQQVDfBY4aWLT3QoG/phQ+kk8WPW6YgAx8Tycak0wkvWQbMRI/d0+ropew8CGEldJ7oxil
Xstavg0wqMsP4h05PAKFCT2uO20u+RLbDLWRArPq+4iOj5Ngp0kDWYzrLZa5TfFJCrbhnvUabD3Z
VAWdd1o1TKM0fyytKXYB/wlC8GvLw1DcV839c7FfuHKFnK9hGEkrlEDhw9lHvvLACXH0tT0rdwXi
3+1ongD3te0k/itDdmKrwqri026SncITOA9GsPV9lOFFNfaMwu5xIk7vJFmDIjooB1tuqoaI57lX
84Os5UyJ7ayzryK6P528ftqJDI/l7siSgDTFY8faO8yX5yPGByEmS5GBqw6emvjUBrHxqvdxvtgL
zIc8UnjXI1gzwBsz6vCtPnrXQg63HV1h3PyVnur1LGIq+ufC4oqmLkBJVB234xZ/mThlMInWOCsc
zt8gXmJf0EIVUBU4gPlKiOiQeP7nnVF8cm2BSPDKy1I1neFCJ+8yO+bVEEWfzYCNDRWDV2Yiu1yH
0t+m8aUTcxPkZxP/HZ7rdY+cqVuMq30qIqHTKHDmlu2/OWDRUjB64cqiLlPzaUcNSujYql7BvcoR
jLRXciGc91zc3QiCXSblKGJsk6BqZuBT2yEYTIaVFMMyjkSKTcyQQv/paOBuYRylS7noSYSYcv3T
vcftbcdvx0gpDsmpcbY3GWXpGHimggOxOYfbR5Me1b1Ychnl/0Xv0qrWRPIB627YU8WeS3Qw9lS7
+R6ycR9m9/X9H+h1N3S2ugyScWX+bKJ+A0Omy6KQG7rQxcImGz+8Xf7JVSYoAL7s8eQboYcD7J4x
V7+icZyOxXXk3iNDK6ma+81L/eUQlU7R4NFMv0J4weQRRwTHtt/uiHia7Z+5du8F02oWJ2X6uVSN
L8puUcJJXGfIXiO+t4l2yDzu+ISygi9c74N9F4a20iAyNdzmsU1AfO581muabQa94ZVY/cW3saXy
r8qM/jAMD+uIC4o1HtZDNvc16Jhj7ZqbKxiCQm5iQGFVZclRI5NS2taWkIwy0UJRf0KHxMIVVORL
sGH3EQnj+36B+NL5WhKB+YxnIIy3wT8gpp9vCg1yA99U+gUsXoaGivkqKKKI7Wv86zcDgjZGG0gh
7uI0yJ6PqlZX8R0dAyfvkjhzn7elM1hJjSVq6HADuVaatduTx7qqco8TbJyMBKb2Vj+l48RYOTM4
GPJR61cN5IQC7qxESh9YydwhEdnnU7kBFe84S3lm+0hcJRG2hRxqdWSnofOHJfwgYULg45iw5Qoz
rGtJ6Efu5QKN9SmeD3754T7KrZjyKWv1BGlwclc0m/ivg9tgKcblTDvAnE/yEZ/aJ9tDVAPWMCvx
VUiStiZMiBVjCR++Ks17pANcLJaMQ/4udpGxhP5hxPXtGDhM/aTRbx2rSMsQ0aY/eQdAguLKB/Pe
kAOh/aiNsYiV9ynGLBZXBqBlwnYHrZqcTAhoqSHFt/5oPu9XlRv1iSmXWUoH/QzfUtGvVc2vCZJa
d0+2eN2k1J+J+LG0NIewnIAGBbQ+wo/4r2DJIoCTXR32vE8+huglm0LkFG43AikMBz3jCCXYS111
gfcwJQzEA/Xxe9e9gSsND60RJl0mawCgey3/50LR1SCSMEpNgcdqVU/2EiCxo5aXPlUqmOFI8mqo
RKl/y83uARAQIvvRoB6sr/oBIwbAbDBFXs46N6D6yRa3EVTik5/f0qgbXxCC43fpXDPqFYwbgmGQ
chYyqUpygBhovsJJYiYxUQH5Z1Eh5fl5A1/M6TpBe4eSxd++N5SPMOkQKS2NgtdXgWzZvpmUvcAD
wItA/PfXAtuikwD3MPG79wJD3yURz57z8hrAlWLFKgKMEwgQzvzpCc6lGabAJTieP6dPf+IL5jYt
1rY/RlTuIOt6Empb3+6tjdLpJPrNt9/sbUHUVTQtdsiZBTTKk0vCIQbtfyKnPpV5XPXj7op2N4HB
wIaC9YG2WYmGa+K1EkzKgj3MCCR5gonC7oB0/8fvfGtOOIF7YrRUlRqrxTpiECriP4O27I9dxHaH
8a/OspJs8QH0UHtn4MNvGber5WS2r3TfrsrrkA2vO14N5EC2juGE67WlRw0FbKY0e1ymMYt4QkyZ
gj3x4SGmHO25YCMjkEDBo/WF5APL18qDd5QTcNEdCjOvd0ZM76mzSXAuFhoSfJpJgawfjURdXgGY
wmQyluB5QoBDL7K8uFEXZxkcJca76KV7IcxE7HCglccw+sd3Z7/zq651xVfOhMrpHtJraxbHqIR9
kKUhytz+EOFBVVHgwLUz650X197dZiIbeKmCn9ECzwGPMbBdEO1YITKU0zeVC67tNf3IkfsvU0wL
TShvt/oBSbx9MI4v/MY3pZhV3998u2gFKLHug1QK39dxrJ53s2EzkYX5skCvsl6LaWLFZ7ZEhUBo
10aW7GA8Jent4XgtChlUtQW+TbilvIY9ht83lpqplnxvdCqAaxM8J1Q8FR1Eu6IvjcC8Akb1QB4X
g2dUMVskR2/asgZ22b5X02keFRcxCqy1YUI9zPusl/dxXP94AoABumxSxxuJBiUzDfV9huh5C1z0
LhsGFMlPpGCInyrQjD58vdP0vBXLIsfth3VKu3+9FPacECHhW4a7s0ZlG8NVh2kIsMeLtOT7vZVd
vn1OL8ckHipsyj/KBbUiFPICgAKEYvRujBPp/AO0avcpACl9KHaoHTBtU6h4yn5pHIC2QQOC5rV+
R41k+4sib2q1oMVSVj+Sv1EgrWRk1ao9nrWIbY/nHuv3LeFRZXfCtviw/wsjc4oMCgEPhvS+4PZU
/sVAu+ecZxGNw14lOYyYWTk+UFrOyw8o9pzq1t2tQPMmsLn4tGEQB53HErc4pJfjoXZUw2mJiyta
y9p9lNsuo6NdfVsEZ587kElJWKCCXJBaKmB8atUA2msrW4/7yFxHhOhi/1P7Xxst+bCAvcwSvQlg
rpi3zC9BQTbxP77F4pJD5peQqScu1t45CpLOf0vHotDoXYSF0TUo+DHczKwRHmpYYSrF5uridIVF
WNpli64rvGFiF/9g2Wz0MIkgD4ax6ZvovfxyuSzVi7q48MpxU8AHCntU6G7c8hnEEmOeypjT0eLg
xlIfeSAwIfczBY7WsDFG1W78FQTMCYBWI1CUiZxW9BVvJZQ+cJyGRctI7MRmSZpK4+bhnixtNXfo
qgR550qx7vQvkDZZwUgfW6Z+eies/A7ICqH/mJXu3fzZJWQ5l7UoUSl/h1vCwaDDu4y7dXJD8Dd/
Q6UKyWjPgTjwMzzZLLxFDtmcbD0mJ18iqlmthk7M4UIZXTJXrgmXBzk/22XReVCWW/acwrqMW8Zn
sZqCHQF5qIvyfn+ATduVBDdEvB8kw1a+zElHFtaKk9J111fNKLd+RksCFgH4BOCuYz+IchKnIw6b
dwywvwJwg+yYmQ/htyY8vvzNGp7UwIEn7xi5b5W6uCcXsyA/nmLimj5SLGlZeDa0brCYhykVgFG6
UNNq3Gb901u7yzqZBwmQuql7qtsDjUae+xemcT8imnZvJ4Th3WeRTFSZsA5E2LZHe09a/OeLsSFi
ZOaWSYSMaXPWHH0PtSUiimza42WEsvnhN7au6QfHlsFaX/RQ5XMBSF9zec4QlFLGoduU9wtu1bTw
C0KLg2M8Ufhw6CnUHkY23VNpI8v7LsIhnR4f5NjlEdBn3sHKaNjMR0P39cgZpZwcWdraZMOxgOAB
kzGvh9gjZr6SXdyFR/8oSpDKgVz30hfaOYjn+EcpHJRS6sTawoMeZoo2tiyio10N5QzzUtCvhO0S
hdlVFoqeVUbxJOEa4ZI4mkKQ3LOv9rQvX9IKWV4p6eK9habsbiOCoTu/qqs+LyePGSEnVzFsC6K3
UqgpsQPpRkriQuEpHbAYh64d5tVxgLLCYhduIHiht2b1550HlcMaLiRwCKT0CXW19nckRweaL8Pk
zy6MkKFrUqj+0PjlLnrG2pi3pnW8umeLTzF+aD1KRQdHfHgDN0d7wgWKXQfM9a4Jni3u5oaJ5o8T
KGkMrIn8jDkxVnfUR/EKmjTtF7s43IXqVdy+NEVMiFwSkZ4P6ANdc1Dj9kVomwNbf5tuTKzUn3kw
Ljw2qmjku3Eki0kRxrG8BkBmMaFRTfZEXJhBGUHYacizVkfS4Cm4si5i0Q6W2WfDt8WwIay1TiiX
EB6DN90Loys7+dHqE4KLLsPBGaWlbUcBo5JSprL90kWTdqiJDNS0Mg6Ro0elpFDehYmgx+psgWi0
3XmgC0OS4wPBUD5CNn5BdU011bFBwKHhdhVjtNANBXpEfM+Ul69MSFYo1+qtyK+hSX4spP1Ljcp3
QRsYlN4rE9EkB1hvl6H+pwMaS2zknLO/B4IaUBzBFoN1l06JEtNzjLvpVoBdJ+eRVJ7V9N2X99Je
KOc8te4cguEAN/XTwTbTYAMntb0igC+Ozv3QZU315EcfbvO93/YutpMJ8jwvtXzDcNm3bjC9/W5q
Wogxw725LYWrfA0n+pUaVB90PBnr5PqpGolQg//I8p2Neb92KA9Ny80tdQVKEDpeFfXgcFVfGV78
l2/kjYlEJ1/Saks/Aqz5R5WpFByymVyssuFtxV0+JeCOFCI0jMdGOTojbgvcTTHk2/5CEbe1muUy
Gt4PtJ2UK6Rh9V3e1C+Pe+1+CPCoQy+PFblhNK2ID9zlFwoqk/AZqNspKXMiPJJGGxCQlsUiwxlm
siwEBkE2EYDYn6SG9fB2pqjP6ebVKz4xlzjMRxjhn9IvKol/kA7CBB4Um/SMhmITM6RfGtg01Ew8
9KPKktYJrxY5PN56NX/97YB+8TmuEPWMp3A31nTa1XhS0HdmD8L+Tk08YpLsz2E+QvpjmI1dsZ20
YfuUydOzUPIhCmPEi9lcLA6FqwfLZKMpGymuo7+pnBonzHXI2zM5hfCvvQls98EKvK8l5mN8xOma
RfHRpbF63nS6KT7ZsUHZrGxk0IOtdenEcYES0M9iEzipvCb/V0v6GbqOQ4I4QnCnE9URgDqPst6h
xOcHD37q8l7duuPY6qxelRfSFxcm6bQ6tqiSBkUjm6rfogci+NlGf3HM8Y1HaPRb+6c/LM/YDnrx
U9h7YGPI5TTMdj66lAMnvn+zOIz0JPMKvlUkMRVq476sM25fAVk/ecPc9XoMXMt814jhbU7ykF4/
WGNIWaFzwpAqFbKG8PI4hCmRUZ4IgqBOHkkN1ZbiOSbB4ZBRdMEX9teIsTIa85A8k/AHjJM3sqo1
lvaC+ikdQzsKBJv0dxZiAu8juYNhmA65VQpoMC+OOjuFfdyl3v/tJqsub+S4mJ8QzyQNapOaZsIl
r/IzETYRmUJ1VPSX5k4/QCVQeQTCyERsgoGZbQ3Ev3K7LeNM8gmWvQ9ZQab28VDwk+PRitEOGJxu
HaOELuQld8p8FgoXa2JFGPQOFVnKmEeFd7slsPJrJf18KqwzlxNnsUI5jRlV0RDIsisKpTyrv42x
00XiHTznQ9cGhqD7USoaTKfB8WFFq2U3LpPe9pPAj24GL6qluI3NyUPyj9+bEcjEO77IRSfLPqz+
Cs5ia+5H9ZZxPwWp9Ib4Y5UA6oqhPdN6JYUdxdZeqUIL+wenvmJWSs1jkQlE7XXHWI65uyQ9lNJl
bKQVIIt60j8xw/mxP/UGpMM1xqblK+LE7M2ZTlE2uibPfdyyKA54Vnk4PDGO33NTtpnQ0eDRl5dV
fswyXdzxVmrjho+w1q4Hl8z2OO2EUQ3jhnBhMhBg4KECFbH74KnUfg98V827q7jwwziBuPxOUGEG
eNNJ6NJgJ1QXnxr3NxA6Iyh25yCEsdpEuYcTyuumRvzfcekrBZJ0q11r67iQhS7EtgeCmk4pSDdT
KBcLQ+9TylG/U3utjWriDCb+uyVsRSEpq6puxHWOfIqdLuTf9ugVuCHIJHeQc7HCVrzZn0+gSZkz
ST68viZrzlQ9U0HyhtZpu1YN4ex1j0znkNV5ag2+ZjAiu/Svu1LG1+N6Bsa1EiSG0f/k7NehCcjJ
u/kH5iDRbPK8IsGKPOwWPamGfVsErYZ05gD9fM1JpeRVC6ZdyZHRcVwOKgG/uGHUSJPLg0nyzQTS
OPUIIUZTkevBYtaVnhs/7v3bdO9vu3pBs10fb3KSOqRHkPCCHattFYm4BW6Mk4xp8c7+lApm+6FL
reLhqQceE9zi7JUHTvKOXl93A5b/T+/KmxCVQdjf+jwK5yd5V2pGPBjfE0x+pFrQYE+AFurTK/JF
M0dkhwBsP6zagF5lZOqVqR4Q9zeeQQI2KZEOdioBzoX4mfEoVyl4P2MrPjrX5/+Kz3ZGx1BFSAHB
848rFl1e3h8Jf9wszNytWZh/3baIC3Ef8GsVBvob7qg1bPIzF8wXG3VKUpTuM4zFddKcFtaybKIy
Ow4frkumF5sAVW0CrB1L7OZ42kXlj4OM17WYGPq6qPjDAWat0g7m9U2WkwB43CNkEAAfGycEqdyk
65u1dJEuGWG0eKv/TG6IMtY56xxzdwW62ztDGUVl7yn96nd/Z3o/fryWZkrSfM7CHFV9KdOYodm6
Z410PV+qen6M6xgweU/1AMufB03b9Iymt+yAvDTrBKTzo0Fgpx7A1iJdyTykKUZhDaj7A/Q42aps
SJI2osudLkN9RhoeyF6ia3E+acmfPkyv4X1blZjj8orrZci0Ilcq3cnIBbuiLzFgn+K8q0lZRZJ4
8v38hnsJHbO485B1OiJl7lC8uwyJNraphMpWyrNrwIE52RIf8iI48FMXA0StKr+om4uDky6/L3bW
oN/iLkwSp1gJqJldBwzQPFQVf4e2QO/AwqBR9sCxdVGPrT0BHoIIqBzP1JQT2FkZ0NdPG0RVnYFo
lQ5mURIb2auEoxnJiCSFPOQlFyzUX7CaBi1w0JFCjPOF8LMs54GhxxnCQrJ/q2pAUTR9r0zDKaug
TPUAFPZVu1SHU+AW7gv4RsVo6bvu4iwPgY6uFrSMtYVx9MQouzSb5YbK5OfhoS+2B9766AFo/Urq
pD03GAPDyWCOdCvLkQ3kSa+/wb5IGaivbe0zJLlQJbaNjC+eVuzKrJK2DqbpuISRwsmMYBKRb/ZU
5KJzTi6bmtIuKPocH+Agp18gzTcCpjaQzqHn5sXGQZ2qq2eVrCD/yeyl6h8Jn/kLhVaaaojFOr3d
1vIP/WDwjjc0ue6ZFv/j3Uy4FZ88mKSBCoYlMsiNXbgHmSxQBkags12DfMSAQ+hLazVGBLKu7guv
rZG7TUSl/78yt4rSWGwI4FUmBk984Zc3CBcZOC/VVppn1vcE/YvrphoX3ulZ87ikETQYnxYCWOpb
b74bU2MwDdYbsavATT8AfQIrOQLVoXZeyBslWIpTrZ/CF0GPCiw4Qq++iJZFkf9KiR046Qqfwj38
JeC1NN5uDVhIt5NqaCkptLuuErTYEVmDY94JaFUSpGSkzdiB6NblRiyriLr7XXEbbshRARORkOYi
yhRUKObhiFwYzwYmFpOZFD8vQ1PxdMIszAKr5TZV9hafpdJ21jEBGPABUdk4FDSCyl5B8XSt65vj
eUs/geY7s7o6dxb26fUv9MzKYpoHT2kzQDQOZukROrYnY9s45PrXouZD7xhbZ4opZEnl6o9gS/+1
/0CJzMvikbHNB4bifwUqMEoKE7rcWTJKzI7NH0BiIAGptDUGxgA7K6+Ph5dLiBEh40lxkJuOvRc2
pEfd8tzE3S4X7Yv69l2txc6rjWWxFfZRv0WPf2oxFm0JFJshxCxZQVz3KZXJ6iazDuJpmWlzowRQ
arMWNrpOe300Ru8h0TGqcEEKjWsSbSHnS8PFUEJZ6x8hbePwk4M8hQYhSTHjfsuPdXKedSy+HYJa
+VjxRh+4AlEO5cWuyhuwU+S0SS7s4NbKAzRJk6hZnkGTgQCh71sfoPheSksERIWAGh1QJXNiqcKD
7g/TkUBO5+PjqQRGqxPN4EsZkjpPUNq3HGQMJT3NPhygFX3XlTsQgtjoOEKV6WdgkSKPoSH/gje8
UH7eInpwnZ8MyERBDsni1ZI/Wv52SlpviAj2ZY++KD0zwLpu0F6b9ffpJe3lXd+vs+tei7Uo14U6
qWzsFTg5wugJhftcAg99mibrt1sO0jdbbCxw3OicsHgBC6+3MEwucJxjLaIZk+Ykm5G0NuJX5FRy
gIPBXoLbuNqxjK3mqm0cNjcxXpukqnxrYrayPYUEI37EIU1STxas/7JyDoCtV5XD9lwrkdYb84Em
/elnicsu6SkLCppAjNyCYFqtEc1IM0eKak2kIYQ4kgezxYoeBJTedfCUdUoLdxmbl65Rd0rDJnd5
Qr3v+pWEGtMzbL7BPJGges3EChoUm0pk84OCIXuOEmsxEGYbucLx2HQ0xJ9OqSK9UPpygXTu72/h
MYjKo8/0kkiFUsuJSkyLYbwRnX4l30ekazoo8WJkw1ChuqjJAyTEajhb8TLCwjmxX8HFIkwkz61g
ZaWnjQN8CmOEM3nwCIiCDUkJhWGYkPQpbw9MUBp8kKoF49ZU2ej9lpd9D+dtT5o0EQ3Xq89XhZxL
Z3Ag0y/BcnQR1rJSnXFW66v05trEUhdjdAPy84fOZlQnqkV4hJ75x5yMqGcujPIoP8aAX+xn2uUE
nz31fcx8yPmYkQ574Zd7l4l9zsHu6+FD7cWFtypkbme3W3Yw9HcxKXAppfPIP7g8vA1NbX8zTzEL
OzcYSWUaUNzcZs/UwNq13aXjPOfIem/oNCFH5pyc0L2J/Ze7BmcLaIEDq7nJNUufFOW97RN5ka5V
D1cxCCisJX8STvql3eafFSjjXMgPAwjbh/VHOw+jgOhNoNAxm8Oc3By+4OnjpceK+uAQkk5hR065
TcLs2SWemZWjNMSWXP/jT3sJKdTq/QokBYBfexpCvOxDlkOuoGThObb2QXWH1HbB667is/cpLjZA
lGqFYpDggcGmtJOiZhYGJlnN+DiaupvFmMDnN7Rpycj+A7SkjM7ix9CBx4WTEf0LOBUE6IilJi5T
JDDBuEkxMWVhJzq5PaDVSgb8UW6ZvOKbyGfGAeJo24SgOC/feKzO5y5+Gpt9wB5IhRtRVvwVs3VR
UfHIafYnu5QVCzSYZz+CHQlWjISk7g88JJUSZ+cSAJLz+OpvcY/SeOcAFUE9kvV1swE0Fp1/S2kx
PMGHbf2riPXG+26GD5G37Ut4vIexCTliz2A53afJd5KEkac4QpgpELxImZSF03f7dYemQyN+Am7K
ftMV98yRo3BjpT1qUS+XNysDhyTywLW14ETTmqmtiTGa+DBLXAQs5h1scmalVI3u/WkdXb234+KT
o1T2YCqvX2hBT1BzAh84+caYe2rdR03TubqXU/LvVDJqLV0H4NsRcTSrJE3Z0feFPd4eGo6pXexU
EU9+JgJ1sDpJLJJ2CjGWGz40cLoU+d2lbQhPR53HidP+tAv79cBgXUNzTQ9kzaaLKBpkVGDBbM91
6YRHF62JRnHsmx+OdR0Tdv4l0bPvqbfJCZu/wlb6lao5i9TKGLXsQxoEuVWbk6bBVh+cTXh/bRhG
VPbfnxHTRGLt+IHR7HK5Lc/2gncb+ZflveTIJ5YMoi46GdLG8QNP6TB9w0A/XiAzMIpTuhG8tDMs
BHJJOFIE1lkL8kcP1r3gDrOgTjdtZSp8/IjyCEVH9sWKuj71bM54arBodA5/Vo4HE+xnsd4ZCyRW
WhqxD5KfE+Cqz8dZ9SVsmOKZtJq6S3jVoHG1t1ONNNpe3Y72HfsWqan4+9c6nzobH53VVGfWQxWx
PC5Ldg17czZngvaSSzP/IddNzzOznpodtivB1UsNTTDEGfV1XLQoTqbr4R7Iq1T3T1GDKV0T4AQg
ySOvwzDKpT2uiWhKPihzezPwHpkhCJ+/SoQ1R65L04RkBtbWXKGjYCkHlHt+0H2MTq6mU39M1KfC
f3ehrKVPgieR3lvIvEaAla8UPgwcSOMG1uidCdhcd1R3eRgQsDv8J1niYpgvB2g+4oeKFE4AlZtT
Slie744wANjLeDKknFG56gwB+iXw6qxK04fZh1tzcL0jZ1s65Hapc09dIQW/VB7XPFP4GHZ4XUCQ
h9i7jDBU9m+FczLyyie2T0U/N3QxKIpBpeXRS6DzxG1ja+ERtMU7sbXb4MACWSc7b0S8NAv9X5Nw
Or7DRa1dxLG2tAKBl3BQNCr4lel6TlKPl0sNA9fVUt1Wg254Wq04c43MKLQ2Avdn4yrM+2eQajTs
rKG6GJgaAYFKGYR9UcOuOXg/GBBYxBJUTcK0pUfaw3VhUb2qg4SDen8u9XobGZ6Ibo/4MAA1zbZ7
tS61URXQyl355BtdNeTX1nvI7ySbXj4DOjoE0eLIeoMteesO5RXkF/zQE0ASSQf9d1zOc0lJ0paA
YojzDAxfAiDh4lqjyXmsYMkfmbesRAT5mCREDwIfQHzotNIoMmM3mSb17Tdy/jxwPYpcx1lvIzpp
kHYZ6HO8Z0a4RY6aFQXtu3rGo1uBeInvIEl4juXF7NZSCmBbYE669BP5wTPRMCRo11oA/3d9+BPM
SAlmUuvVXL1PIgdcvNXITXsHLzqMWdlDg6acMXVP45TeO1rzXFQiMJgcZ0V5Nj14wKRovEdYRt5q
/0lQkzxkuIPHWMWQHSWViSsG4rZ2/TljL6azK6RSJEWCvAcfWbtE4FlfaVAJEdgc4PoZqwvMt4+D
+Zfw9vglnX/3/PIZNMinVPuYHGARwHtAhxqtmvwg7NFJazUGO81tjEqUprys9GposDNOMOO/RMqT
PhpaMgZlCfovpN9GvulxEWVcFdRBG2gT+rtSn/HT52XOQ4ZtrpdmVkb2rBT2p5cflUgi0m09z+cl
BCjLedMwXWBqbzwhPa+05p6HQTB9eMnjjZsbfm08wd1lTQ5hivL+xxUT90EruZ96TthxTYmG1GfO
/Z7URO95qnRb7edDbNHoX/UL69zVMWhLJrcLWRpm8zIvVobZmR5mDi8uUqlN5NhSm4zmJtTt5Zjt
fyt6ekBd4sW4xkzJAlWNxBhhcg7EE7QrMGeZS9j9IuCTdYp691yE/wWhQDVhky2FJz1SHjXlvDl6
s455Ng+vQz4WYUAJs4bV1qE4lh6mthtQRQbcfV7Xi/aaQt86sEan7cDJsiZQkw3iqenSGyycfpHo
+b0wVDQzlqa4QwdHlNYqOHE5eSM9hv4k4PZ0zte/bZ/8gZLpC/YUNYyYCMp5ve5A9x+6crc611Iu
AcwhxiNj9vpFskCy4yLzPYhSc0oxJLVzsTFPim9qU++N9EPxCwCyAsQTyKlpWgOZ+NG6iRYvZVSm
u0+tp3aH9KK6w4s9hihZa++dF3zf/i+DXQ/U/gTK/okMbMSleDd9DXtEOIu792hbiNxsQkLpFQXu
epVY6ry4dwp8aj5ixM4PnkOJZbtVaA5FZRgrwFpuFmEZzmYczVOK0w/qUbxz9V6GjthVPbAKRCeF
c+fOrISVZEods991MC1qME5Ll7wwwez55BvucNxKdEPhYMdAZfKB2B7gk5LzTFyNhy1f6HHfegkv
W26Xqijsn3oVF1PKgSrwvKGzEDFzvkbGLXjRx/cNMjauIaipwFg/8LDLFrCPeculY6W/A/q1u6Fa
gK82JqAR1R+mLxntw1uUS22qjEQakiYfSz/nIhfE5dnDH+yUpc2PYZ+wm1vZ3+fGGJD/8mh1NVOj
x/npQk3fte/pTjjX9E3Yjg168bJyLVcUqPNDQzDUGkfQ+btqrl99SbYPy4Jq60JPuh4omsMr4rsi
BGYlCGxnnZpTRXt3PlOviH0dR5Z5STIwyiSPVJTuHrkyiBhxHVuZ7XU+2iv99qElIlqFMlQ05hLu
rQbEb4nhuE+VIko4Al+xulQWxJy5cjGQZwreAct534llBJ7bIsewyFWlrxyE/LUgzHzxVG+0SRwW
riZ7quoV4Qh9sPIeklM3WPOXTifw+gfzAqiNPLejKL1rtt3y48zSpJQqbraAT5lnR0BCXdzPVOMF
O0HNo3TSwyM56MSw6a8bZTed/+BIwMcxq7ioKPcrwJAKl+2lfjV685tn85tC44/7Z8S3FKRPYfkd
ktH5uF4KohsPdKJwSYvd0GTujN0paULclkeWd4PJsKBPxB57CbiAQx6g4P8IMzqGftmEdR60GK5E
aX4R5mETYR3CGswJU40I2+/u2SFci/QxLvNKiNV7nrG6D6GoT1yJkW7fC+rOjkejvM9Xe7vxt4Ne
JOEVrwogQj3q3wyYUqOS+dfDl4KbdARHoOYrHc5Oj/dQh0EST+mjphO8IQwR1CkkPN2dRTUqHE5V
Tk3K5SVVWWyHHoui+yHSfjoDMrTN0GAFNfLYhfcsBGjuHAiBWIJjyAACh8aBNud03CNeESpTS8vE
MhAxBLN/1XAOhBpqQoE+L0ieLn8gmS9R7zi3v4njoH3kis5ANiXBzL8vLDrMlUrCIi+09K++vh0i
Ow7RcJfSM/dVU4FR6LZ6lf0jtvaS9+xAqKhuSc1d+2LhAa0KwThfr8KQ8AXARDT1EKkTl1BT5III
ckS4Sa4eG3HJdYPvFo4LN9GldfAYDeNI9JFj4SE1GLmp5aPhEP/eEBzqWaYdOE5bJQ/iiUnI4uGF
UlFEa4neGbaO+NU3azw7TK7+gF7BdRsGGwRBCOtduaZ8xlbHf7AiptAJm+xD2MCA36XnWoXrOXd2
reKk4poCKx/WL02YR3qmzBTRGlHLssEnLM1URFniifRlhE+R2qA4mdOL4/CvEC1EnqFEY4FH+ddZ
vCMOXChoosLk+S96iSMEOzEa/BygV3M8Hdf1RBzXAQWvW9bEol04Pw7gabld+wi6qGmLg3i0E08e
xoOhjuOHJjd4MrZUVjAmQuTy7BjWYW5cPDdqUGhjlSoLBQayVl2RTwTi6RRPk7+ifz3tlY7vsBQU
d+CcDl3zijzA2lfPbmq0TOZakOuObBMlQTuN7Z9MAby2Kkzs1qVwSlOcrC/6FTD46fQUh7K6NtI8
DT+KOy43oVrkQoKgjpTWM+R4stM0dFmsCZGBFlVowKN8nBIYLbAT+NhYz/TaIQTsUx+UCyhnQDOx
Aay5E/zn9WWUJ1mXAIMTmZAszwbrwrSJQqbS0gCrLaEPhm24vGB4S/kDZqBsTZLapBjUS+6Wrfow
h6IaFhSpKwiC7+XT1bmj5jwRKcyTx+Bel4Tupdj5tlbUTKYG5EYi5088z1eUg87j2IuGv9HLBLLo
DXQa0sxUQbJ6Azhw2tpBSAs+Pm6KVNlEIb9d85h0YvXhoXI7pviGbm32nfI335vSujso5DxZq3pX
Tro1PxfRaMF3Cx2BNOeq496dILh6N+O/J0gTNeBGh/joDO90jViIOJRChzjDAvuCfHJgZiLQANpp
CQ6uwbu9surwlf6658oFwhQh0gbNPG58EDRGxCh93EBvK824nRZvkD1UR8S3mbNqxRGXiixAYEf6
DSlfezyGw5lBWJ7qk2WlqluB7FKzFa0At9GO1NfyjEaJM3OR4vm2l6pWOz9YxMuK3/PHOOj9iDcG
gE5ZfGJKzKcCliquNCAIv2W0TSMuqQeKbiv9MQlBJSHZEot77jSjuAdNOFvz6kCbJQXxo/NLWyoM
jMd7gjz1IAB5tKTd/5d+C0aEaMiARHEKoqMNHAIpsxvytRuNsVA6uBn+EqPRS4pA0NZVu7msfKpF
HcX/75V6DD3up1Uji3Q7WV3u0rl55BgQkdyPy2MJA+lZBPMs17waRJvZzWall3V0Th6PKf3kwbEO
JF4X74oY7BB0omqlEZiRjnd2Pxqr7+TDdS6JwdgFvxFIMAEDV3ERmZXL5lC1XbrUsIRVz7cCkko4
YX1t13s9s6+97ZPQQgCYDWQ76Y56562P3Qc+mH7D+uNZoT7YQWNy32qL6Go4OkeuFb95WNR/CznW
a+HtP2LBlebza2XBLruMblKk3LMGPbC7rbB2/YatAV2/NlHnDpdS5ZAUVN0dBvsqtOLZXWNb7lZT
txZ1rA6o8DMLNmqsJH2EWUwZy0Ikl5mnF2gZEHsBnf4R3K4daNTNoBYG2d75bFIl1YIbWxDweDYE
g3D12puvgjtDtCB/AI3BOAu24+aWdTfvgdtXv3m6qigjoKh9s+4Zqc99+TL+Y5fmsu4LBdpP6pPP
uUZYIk4D4M3NpC6Uk352DC3gLzFodlIMaLnTZR/tPGLYIAIDWkioq8QfQWO5+28yfIfd0OmFO9xZ
irNPxJLl3J/Ur3VmoDyUk60RwYIhwhGtXyY7jwMb+ttKv5jwXkPOViVrQZXWh4SEZ6ZL9+Fp6VK/
e/mCmnj5kSSpm2zrj+bQaHeYC7hz/e+SrI91kJpqb35Wber62n82Gwuqd1zqmF5GsjLiAmzLiiiU
1WiiBTXzfbIdnW/P7iGIG6wmyNzG1h0WRX7ziOABqBWRFS0G9/DosMbbRLx9+dGA8unke1KURQBz
E8oXNbFhuMnFK8gcI7pw+HZx54yJD9ACEu7ATTPyOoSUE0KT7zgJcw10kg5XnI61PL9f+oWKuxUZ
3g4jVs10XpRNn36Ifvogl6NA91mS7B45nMEhG0NnB1zSa0ejbzoI4n50hRfL9ZRYSYArluL+mnig
28jjEcQmGi4wIU7n/kcr8bSPq61oqdoN35uKO7grtZuvAUgm8b7+YcGKj3YIFafYqHb3FJKasuf6
SzCT3xrL1qnfGQvBWxaBOhT+qlaaLj7S/Yp9up/OILJN+pY2+1Zx39oZQoRNUeXPFAXMhnjiEEGM
9OUQeKe+KwD1ptXxmqYWs85AhxnAhrpWPxrrws+cqNruWOzbxgmDbBM4ZT2YdLJKmhufosqwCdp1
yHyYGL/eTFhVj+N7UsAKolGrepkPPj1MPxBspD3W80wgQwQ4FQbpQdD1t7gNe8eql9bsMfRKmCGF
omDZ6pvVyAGGZ9pU/gla7uNkKkqRxvcyB7y2ItoH7BN0DES9KEqI4HWq/Z4m5cg0SYGET3AIr/Gl
7r/6wBzbHTepGgL8DH0rfeCsp1CDpo/WXfy8xyUkp3e1lN6vbejn1yaPEOt8jrtaEzDYFa28mNqy
UUwi7T7ImlKmT8SAryCaIE6WXsUQ36zaYpgK9kdZqCUMghPO9Uud+Bq8WveDrTfn4kmxnluj3zbv
4lsmQiTvQ8V8UiZ4kPf2p70lkG0kxotAv/wtWx2aMlze933w3SdLhhkToXdhbCtWJAQsFXk6Unuj
R9FY67XdBvvRmag6/Hla+3YrfJ++4LxDUuEBR7WvS/DjbPi+y0/3Imws98n98wRdUHGkF2qWpXq/
lCXu7r+wg7xdkiPchqhlsHmoy2QhPvf6BP24YQFsdcIf9URe7E9cUwIhtU8c+qbWF5/J+ZhthYWA
TqpUydoRFCig45BCv1uFIPSLHpo3EallgOA/jkLDOo6uLwNNhTfuO1TCh6QPPAWkbTxjLzZhTg8q
sG4gn8EO0/mRrdSD82D3HTF4psUiZdVyGj3R3uhHz76uEibBQfWvZreHTXJflL2hnrliFEi3cibD
I9VUT4dl5jR6T2St07KVKPUplq5UsbqNW2sXHKbhueTTrNXZVYUYDhdW9zRlAyVYTbtI9tgnCZ8w
g9+Gup2QNVA10RflpaZ47SELatIf+bPfBvAvpswc+gwocVIuIPpAs7UmVrcIXY7AtqD5RQvgTei+
0425c7wWwSOncY0zlPNPO6bmgxTqhJL+HwZEvWPjO49SFIK/BODomcXLiSYdQf63t7cGXBhXorBQ
s/TKKE9eZhPMAfDwXgOxxSaFLeR3d53DwbhoiDMTE2ZA59i34RUVcWY3f3kSO6ndbTjyWzTr627K
PXKbx0MPNtAa1e6gf5dPk5p93aqT7rG247xqY33F7D1f0ZBEs0j5exSG0A1DzJFIa/HAQTiR7GsJ
quWgFGVVSSCbPbEuN5YvA8vXewRgaixsj+FKuGKlDUHssZnC1IeTN8fM51Nz2lnkoSvJM5NSPsjS
i/jAFK/jNbW2jKoe9uS9k5+ey+/LTUGCNcAg6rYoJ8g7v+QpezDXkwKDWJPQ8OWj/DqNOA/oXgfP
StV5Jd+ejiQEaJMBD44wSSdwTZXPZ7Lfv4po/YRpDg7ju2eO5R6FPiEU2r/KX7TNEXJ5JBYEY/3x
gi41PcJSqriKVjFMgtu4ZGCLVbXK4pAoNrIETlwVkqzXPYBiYZQiGn8cMvkwTZHd7u9YC5dUAIFH
WYAWMvMI81Kk6ssklPFy8IhzeCfrFlqyYbUB2W5RYJCYjzGxHIaZ82t0Fo0rjIkHrW2lL9otQ1Xi
Eoyr58KVtAro7/cFq9ld03bo+E9NJ9jmB+utL4GssL4HtMFtU5kkjKkmH4vFSZ7FezcRt02y0s1r
hPOzQz7j+/bvpwck9QkGYZCp/MgNn3KHrZDtshMbq4nT/+CHEvNNmC8DF8rGDwV2loe7YQXBvZRu
osbVcW2TcBbgAKoHEcc8t5qQ3icyqIfuAiYKpEApeNDdI6GfzOwjOEiGg1ufwSEeQ3gH0N+NfnFE
WPFranbwxm7PXI8/uTNbeS8SLvA2Xlw8XsxVSo99ecjSZ7HudLzFmaDCwGFWO3dqe/IP5tTKrB5i
HEWpHRbX0AJLIHNLiz1v6DE/W15j9neXqIAKRsBDwZZ9zvaHhmOsIjwzc8rL108SJUfbH/rjqMY5
14h94jAHUgVQ3m5ryNghCEvC6XPeEtuSTmNnlRIF7pSh7xLNo3jmUuO/86eI9B6SgLoQwW9POdpj
5/xwWFDBozq6JcNCIT90AJjXWqZ21MdtE5JyuJg71hQT70gI9b7iXuHDuxYweP6TpBY2pD6yAzsM
uB90PD/yj6PlSM2wb/FnvpXkX6ReUe//p/84YFh4zBv6JAT6tOcOwpaimDBog3YP+NRbQzfl1IjD
reGu0y8aajMKkTzhrjRfveCReBJ94cjfh2+lIHq/F2OEdo5uiNxPfV4KwB1S3uBBHMbvWK9g4ZYn
LVIF9KmEFGeXMwnK3334g9RjHu/7fuTHV1rvvqoeQTpBgkxBWb0Pk6Rt1v1p4vMLYKL1Sfbz+CYx
mG1TkA5g5pkXuvWHlSSMoByfdPWPVd/A/rIgeMqOaVr0bHvqfQaN+hfgDKfzkC82UR1htyPrEyyK
FU2FYxECov9Vd67AITCESPrWNICyILeTEjUHDvwDgyLIM3qrSLbYnJUFi+3IfT2QFjNTzJ9WXdu6
Q/XRq9Oq0rGu0BYfbBB2doont6Lt4SsUb33gKqNFEcUnabALUdNgUUxORHWIZINPkz03o8fwxN/q
YSBBTl51c7f1zIfnHORdRuVxxF+Wn2SX3FdoYe/yyLqMw+qflqD3Mffkt+YzuCd2aPPbTARcZkuT
RY/SncUH6kvupcr3cjMIYtzgHVChFWLCeGy0LI64PBwhR89mo5pG+McOHkOYVW4xCHt/D7RSR3HG
FvYXf/2JqqnDrhdpmTGpoFGQY+mvtfa8hLkGsCRPol/3Hkw0L2LxxRWxpzu0Sd+qM7Lw/KgkeSgl
bk/ln6df2GhKPsqJDbqqNnPzgEf1eH8K4ElL4W+RS5yGP3F+WNi5gpppzj6Y98MCP+xf/HHNX19q
1E3CPsmh+4BHtW80TODb+75M0JtZQxi5j7//fbH32s07IjNijHai6snq136a2MnA686E/D5mbCr6
qzVFoD3wmuiG4RorRXbsBSPw+4J3yTkBX6xVk4zOvNmvq6n7kqyJVvQB6mLsLAG6IPOU78d6JKtm
6yS6WxTF2blgbFmkiGE9wj3A9Gw0pUbv91xWNZ3k1jlIoyO78Gbyt7wDZ46v5gSbRgoT2wcOa4A5
xK6BpOQxJH7fK8KJZ0bbxlaiWKvqTBSMy2ysp3/QEffWj3hayj9gIRvbT4jMHJ9BvYZHtV6xrgNA
m8eeKfpsUjr4GhxT3r/khpxn6n8o6TWwWXwjUDx72LNait8fZMIqAtUck4X1cXnLX6nYFrSjS2d4
YdvuH55v5HxhmAXUN+9S9SZn/AyKa/LHCvIpdXNtPVXwBjhEwr/qbh5p46FJAOWkCued5WZI5d1V
qXZXyg91ItdfgEsdXAnPmsMJFg8/8Mph3vZ9kqN6MycxDDcffLwuezrV+7N5KXGI4nJniRb7iuq+
QsHeV0QC5kIY+1EQwn4RK+j1j+Bm2kJ4gg0rjp6F1fY5IiYp9+YmOLmVAegX/i+1NJEzTcML/alV
MW1S13Gb1ALCH8CduxUT61ijD4iS7nmqjCp5uOiAgvrTvcgupKjdPS66v7xSrpsXI7OS0cFN0Uyi
t2dD9GlPU52Rw+TSSD1uVpMHi/U7H7PbE4M36m3OGzKc7wQuTG7k0f3KFhRfFAhagwW2JrrbczqD
WDVd6gkqJjfGNCo3R3xHoYwq+0EpcO6YB4jmzGMwclk9+AOOYWO/VX9giSrUkyHChxy6rmx8MwS8
EoexvgVwcXh+Lt9+QPgtTa6ZlqLtlN+dVLLdlVpcf4Prsff0r7q4ea+frL+A6AyflqllkVo+7DWL
wnIexAtLIeWvSBk4vL8iXY8MHj52O1TDJU/5laW3T0Lbwn74ziAOaYKhnAxmpg+QR3ZVD9YKtU/x
yQQMwOx9rMw8VoSd8+pElQnktiS61HcPeXVAL6FQXs1OWp4asosGVUPh6Ong4AQW2UbgA0bIfj62
SqtWgECaqeJa+EmwWWTNU0G/1dDmlJ5qTFeHZ6HtG9KPBpS/dhQheVeT48Hib6TLnADyXyIFGuPH
kp0skc5JLniE2slPMxpdjskBPsEogIQswzSIuvglgp0APias/7JcCNNWrQt1E+ELGsYxN1oJyFwm
nZGzRybOvQGO12l21Fqd6vrnWf4YKjyYEis1kqo3iwJxHoZbKnweNsa0YPdzlJhaon4NqR2nrY2x
l8FI/kJRu+37P8iFpHxsfbtB93uy3MMrVVXVVR5p6El0LDak3NmMQ3nMu0PayOOs9qWrlBhWBRrE
+9Sto+ImITCCrl9hF5ioUO2p/ousxG772pQS3f6CWQFJVuEpoUGnFlbXsjBB04UEt5YuMPoK/eMv
RHox8HayYjrZ/1n8v7w8jnT070YhurqMTmMa1zBBkw4Tjah9fT10vh+2HDVvyryIA+NZQ2TrzSak
7e7LKWL4Z97t39BruJnvmTcDJHqorI5s1xIhrisrZn46fc4q6ij+YRMBCY4tnFujT53zogWZI6cD
aLrvLJJlkN838bTYP/mo1GpPnBCIl31Zzmj9N9T5PsejR14Rw/Z/3MAcv2SJG8BvF9rAxf1YCFki
7bStWpoBwePoIchLaqojjGdCExq7Rw7TKSAfBLK92WFQb37an/nUaN6UAVE415wN8w35waS/iR05
Qmv0kWnDZmgEFwynzNzYqh35aKIogJ346wci9pYr3W4eV+elUk9MuBxauwJ182S/Tm6yV7mafj63
97cPpVCCIafZg/qGEtLNbowMA1BQ3qO8h0GLJvTIucgsuXK8YMdlUBIywmaQVYM7PQJKreb88v+j
5fOUXn6TjlJXQK56oQxMSfwkDk0nAmAgrCZtdmGz/Gu41PZUL0yQUFJmN3GzHKe+gggTv9lHqu9y
H58F924uhWINXqgog23kQGRIL1ISmakgHxOmGtqaRV3XyXY4jaeQJ3GpQwsW55R1zAH7rGx/OgeW
JeHueXYZraIJ4it9fYQxeS9bBhe4E7LusUoSekM0YisbfmgNMcb20ztrIu5v23fdi3YiDG0E1N7K
sQ7HBWTFXwWudfn19Mw9TX+jVKo67+aMr6vWU54imeJK9wlpqUy/63NI9OQx46kiZkhROSPZHGkQ
g40fE7FYRLN5uEzMcS8Guv8FjyEoLCewHiW6SHP3F1cedoDqiUrKdl2paZ5uEIryk976ikXnhZST
5S31phwjWZ/FvVoQBnuQloP4wBxeQg22RmVmxSFKxf93O94/KGmgnIoMGzm5qiUVZ6Q2uBPJ9Hqx
1NuYynKfBUaBYoJYX/0yU5GzQWw4utgMUcylm4PVtEgNAbBbIL7/L8XNPI/l6v5k1FRXrzwCw36K
SdI5LWiOoI1Fpyw5aD8Uv+Yct1oul8WJKdMIoKR3Yx2JIhUOKdu4eNDlJwwBkddth8O6gTrnYkOi
msnblclfMrDbLCHT91FczwOjPvy0yJZ+hQqLck2IntlJS0QT/31CUB+L5bmIqZLwyGMoh0F35ktp
YjmxQBZibOYONtAU6utesRl/AoZqBRhy6vgyE1beoBy6g8nJLYH2kOIp0CORfLGABGdxqQzFY+kS
r11p3vZRBtj90g8I0bpFZhsYjACdfaQiKmAMwFTZAxBP38YW8WMFfu6SsNokX7jqO9dfuakh+ToU
iFs2UtgWx3ZRbVzFtVnFv+2rsZMMCgCrIZsVgmd+YIy0a8G5n6VmHY22wS7mcTcNmlPrp0HiqrD3
vPfZupOyEX04wiJFB3DwuKJx9kayP8ya3Yw3Wfy/3lQ7YhIOrhhjo+Zq3ZqQ9OjqAXk/s2RHMVyL
5lrUtjzstD6DAyGJ/5rJ+tSF2fxfIrbC0m3hO5EgZZeS9zGo3eQd+2LPifoqLif11kKQ7BgCykxj
ZXhekCbExg/QZlqfo78Ih54VAmcrTTy6+x+i1quKbkYAxASDrDW5xA9MgUy/CvTdJWaiItgji3MZ
LzBOq7OzrLIy256IjDJKdXCIG/ptYJAnjZ0Rp6UmWH2vev4DDy0gC+23Xp9GJXrtA/uAo6i01hga
8r8ei7Hb2AbNS29rBQHzvz4hOscUhV6fA0G4f7/IzA0HEW+05pOsRuymuy9fNANTBOHy1IGfsda5
JZpA3eWQt2glmMTiPWbPsWaHBs0u446QWgwRUf3OgZFCp68ZxdlIFT4OuQ3lRrKpNE1N/EB34kwE
NwLY2LrBYXRJJnbFtyX0IIJW3w9FwMwTaiz2TZjOYySdPeWBOCCuY9V6ddf/7wfRVuDhAe8rAjhy
LzxRjKYIaIk0BN+yspCAi7kkSSxx1qqM3vxvWE8Om/j21NnU3bS1b18+4MdYK3ckGXlWE4VftSXf
AgoNM/bkH9rONzrSr0Rk4ZPrmJ3ulCdTo/41GAjp1u1pKGDjVHQH5Jip8L8XchxCBoG2+Rmlpio7
uLxXVL5wDj47sFWvovavAll5Sfgn4NYojci7AzZ5W5KupcQQ7F6wgs3zfF7188u5ruexnCSFZfVM
bYIKl4Y4guXFc8HRXovEG7Tgv5FDYNbnATXQqvtNZETjba7jq6IIjXs+rkhk6CTJPi9PxISw1B1G
ksHbADdfgdrM5MWsdV9GFAfvBW4Ns7kJvmLn+MzwcG7AMx0ZeM6s0HMUAyeZCaOntxm7vdmLJK76
8Erx+Kd4bVDiJavAApaad9ZXo96O31LH/B+cEZMrCJCYzrxFVQY1cRj/PVXEgcwaRcDK357FRwu/
39A9UO/la/MZrOF0tbHqveU+eD+p/m1/QKxqsmJiOGj05zN32HJuhcaqNkvDBrYdmHszY3hQUMwm
bdfI6MhZmp6HKFDx6+Yx5tt2LG0URbnLZqHJNGGRjWwhHPDcjHw7Me/FmDu59aCRRemNAKkn/ei5
AKIHdEhyLx7TN+8lD+psDhKAB1cgRvk/ziw9VMnuZ12C2iJnGYKfjE//5ezNGaeUnUqAc8KisGWA
AH3kjhPqkGpC5fX/3Qx4ZlnihDtlL2JrdzWJsm3yUK9Suw6BXCFQ/eKvR2iUVO/quOB+4ReXh5Md
p2oMQHGs9jbtSN5T5VgdGcBCM739cWtqiTzcJ70ibjmbgYAbtXQAwVpuNynJx2o4gG2V7QlLYRoM
ga9T+W6KfLYctn0SeJ1nputBbEF8IgwnrU42QoZZT8JPmwmn7d697V4aZ7JtPUkC4PZlWplHqHFn
HDVeFSBeJIja3+WX/rL3kZvH82/JQbzrrmVqy8ACx+nIYsUSgzj86HvQxCZHvt11LtXZTCe9MCNB
IcGBqhHXY5EhUwp6eGN9633iTrr8eNBsImjRFCAzmKljPaRRYVwHpN/eTpyLF/LK+N+Y927YWmHe
7k4gVJrc+kHpusxvoD8iADmECL/pl13gbQbQHx0nMYDrezCJOaLlSCcFtCPKh04G7+2QdswVuV74
/qeUoHZy9LeWhcPCakBWgU0X9bqekmvuaUXsvmWC4JQr3QsDDYpdeFYLn7k1/b46fo+vC9RqRal1
fTzxd5nTKKu8QBBIky093On6ka5ozNNer+YwUtNNoATdr/rMg0hqhOhNWTuNO67EifbxYx1mTD0e
WhhC27BP5tfVz2f+oYusYsdgcfm0P4ATE3miAxv6f+qoWRG2Al27mQyJNJmoIxSiqDMuzLP5Pshz
K8FP7R7aBPziZzBXzdaCHXgGgsOVXNFqndY0KoZtk9x8IvXAAvlwFhBTWD/PHpICRLwMULRNDwZI
UFqEMc+d9T2+HHuxUjPimjSIIkCLc/do+qo7o0nGds59EzqnoLkp14jJs6y/wPDS8A85sO/Usmhq
Hi129Mqe4I34/Vv8UPeyF8FAzxG54IHnINZ7lEfDsMEwxydP9CCBuMYEnCWAkJe3iWfpKHcN2uwm
wykfKlWkKgqhZS1oiP0dbVIaIN5tgGlSHDB2Qg4lQgLLMhtbkH8hQiioWvYGf2TTYmXn8S158KLD
6Xs2YEkW5qr7dBjOdROb/PNzyh9p8yiQpnMNau3GWuYtiDskJMylE1Hivifd4omxu2pqw6KWh8uu
1m/W9sX7BBr0tVzOHO/F/JbXem4EpH7S4poJ7fS/1rmGDgxIS9G3Q+TDI/11pcSZWHrME7ALVEa0
4nzB+EkjS8OV7sgU8GN3vrb6fRIr5o3LAndgYnoWM6zZ5/YgnXfBKYQ1yNT4sL2i35/dVEZzWrlP
3vyEr60AHFb45vXpj1B6g63zMBry6M9b2C2WXzCUgPc5BM+K+F3HBsrVWjeiKcL7BjyLffNJmOkk
r429j+xWElYxKueGBv+inPs3P2xTeIZBI3NtOWvkg9QbmrDd56kV8j76H4pwlTy1Hfv+LLuGie9t
1LakK/xSU2KPxzUHuiPnxUoMpuZktEdhCokMPi5EZ0mxS+Tgi0LryxsMaOoSWAwAdoc+sKjLUdQm
3baGwod3Qyr+6B09H4a28KzTouTnwVErvOYiEfOfYv+QLrO7Qo2l1l5iof/0F0xZpl1s1pNOLAZq
ZpoJ4LUB+x+CwMI5t5HYRtHJnvDd9vJ34D4YRnxtiBw05yBB1orJvXVlXnuAtzkIkSuNwI3kAklk
K5iJq9R5Fv2SyZldoTETtr56bWgpdKllF8d9pMRLd/Wwp2WztyR66JhhAqU1qT6tTft8dFRSDMvI
EYCCicFySWOCezSnl1ifjvssYw8DZQxIOJe6/M7Ui05rJFQ1/u/zybLgQFFqOjGJItPyTcD96meJ
Fk2wv9tCMjfHDvCNXHnqzlRp4PabPRBLloupEn0WhkjHBboHPXgqULk37IiC7AfaUtjLtMhE5DU8
Tanc+5xqtrAr+EKqjzbX9FuL9lIjJUBtrFl4mMf84PkVauOM9A9QkTUnbF6XMwIetjm1+jw2ehY2
iT3LcYGu5mSLEmQzoAI4stLXfjfFa5xAGwEzBCrxkC/Ip4cfUGcGNYAOVFvkiwdHAtda6W3NfBcY
0FSGX2aZbEUicvnK4EooSFvF2uHN8OmeALWmKC9IdeQHIQYZjL92cafYlbOmDUar/lr5YF2dq0mH
o8XSypFnFruMAWqOlEhyWpSZfYwUaneRGL2Q0W2SuUkGCPqQFUDw/n56gs+I5qRS7I6EZG0QdwQb
DYJuU+V8SZ2dzvXQjqev8sjmHh3Z2U7PuxhlWH0hCBgM87thwqBR+Yei5fk6bu1XZEcOqK+/wE9D
3JHZ80E0oITFkl/KX7Fy0YwHzx7zvHKmTgmJRL3BaPg/ZMduRiZjE9K9EjSdBNlX++E86nU5qBYN
yfWPJLdU/apTpEuVxNMdjodiB+rpYOWbA4dJNy6h6Ce/Rx/rtnjryst35rtyIcCYfgijRq6x2OZR
pHvSQgJAYRS540Jq7R+8y8EBj3xJEEVeVVB+xTrKMdv4tIVhF3V+bM4LhN4t8JWlmtUy9XfgG1E8
5YI+lz3kvB+Kb6GQGkY0kLrJNO4njHifw9r/sZMc2ORYQ5YmC9XWUa83+0NyFnEgZB7cBjvmEf8t
AfJDLDFnwIaeviWdL/FDks5BIpc0nsC0zA2CJCHM0iO/PHDz6xF9dxiFDj6EOq2VNJSCCBtdljVk
kMCXg7hW16XHXAeiwetuXd0zu5kBrfVqfVemU3NN6+d5M1uzAFme6xOHchNSm1TgtdzuOLEodKfj
eKQpK04Y1TonPx3DBkc8+ASXYV5YOSMFOUhSIfItb00Tc22FUfKomuit30z7MRTeuNRmLQs8i2xi
p7/pIZKb1JBuTdFVhiaNq3DlvbDE29DuXrrtDonwHGg2+CUfWr0tzd+5XA7aRTfX0dfdB5CRh8bE
aCqL31wftx8OavSvkIxq2V1BBoMaO8XzEKg547efC3UqQxIdAUxcB4UUBpXQnSRxerxhL6F6jwC8
MQadgoXqoFkx0yaeOFJa6YdGsXZq3t2Yg2fUEXcztRk+nloHP8O/YZO2cCO4xDYSQcJaGf9kpPOf
WidtpfSMsbJaEDiMGTtPwpHXG8d79xuwGraR82hPMopARHpI7By3AjxrjlIFMSMnG8HNZSLrQqYC
UCATni9JjGJm318DfyJvqsfv8X/MNgDnqxed1ofpvQ0/93t74n6JeUW39pbEoKMAQ5ryV3HytmHy
zgB1QoM2nxoiNlW/6wP5OCuuPfY19gYTCMGCTjrv4Q/Z0rhm6AFl5xEXQRFi27n2KhiNcmKW71dW
rDyKj8u8AH0/kOoK9hN19PFcj6DwT3AyHrP6xAk7v/BqnpEKixVUhkxIDaR4b6jH2zuaK2TNjeDk
n2Ny5a7zXi2HSSeQRzL8/vhyqH0YaVExKJnmKkWIoRwgVXZjDayY8SaKygYkyzu10XOQQuAZbW3h
OJ1pWM296oNBMqB/JD4y6R58Y1t9OKbqV+xyHY57QjCsg19aVybG4AIk5vu5t3UB3kJsglpYMckY
vfmDpNN5SRNQKNix0LVs/8Rgf3QRaZ7msNcdqpsXG5Hhgq7pSlVJCk7E+q4llIiMh7QO/4+sVEbm
vRpf7YqgdC250CVA8E40olUbSBQgrPDkucPiB5ykYFyFVnfsHLMZ5D5zxrCbjAxrmbjS+pxFeWXY
yiAXjd9hfpEcFCLlGCqAuy+G/J11YpOWbY8CegK7PvqtYx/0OlZv1JeCekKuuwT0ZEnkiioNPkAS
n7RFGgRryuT4g6pM+i8+yeC+j7qZyCRdQqL/EPEY1KfXINKM4wL5sopKqktO+aoVPkDYDWsIomSP
PnEBaqATAQp5XDfJUBu6W/leF1tmPNfXHRQdzC4BSfvB2810kMW/e1Qk+GyDYVo3u3/XImglAiV6
6RI4DflbGhmYxwf7oktsTGDfZYOvtB03O7F+fY4uoBUrvD5vIrTgo6Wc1qmggOJLYnQ2nKPL/RvV
yBxVUN5oejz9ghlEV62bEHL6NyTYQjqEOPuhvTQljP77R5NJq2WDA9+nkWTMGg5ACEIw6A0dwXli
354VsZl6TSkZ6OqVBPVFStGScwka4yGPHLi5ks5llGWXrTnxL1ipdQD0/gJTA1FDkWgLRvJ2fku4
UcvZm28g7sijQ5Qo5IcsS9YsZdzPW14N1yxAHg/7cylFmWoFh292+f+H9fLbKI34dUUfTYh0yZjX
q5oGgMjZNN5I2Zb/KyDMZ7An9M+PIZzv1umC860O1uF4bzyJW7jVOTs5xqokIBfjlL6w8EPEW2Il
XkGcXXOVD/jXnqDcjgu0fArSC2wobE4hsWfD18G3YBOjCqz4H5bP4oRkuoU9z4/p7cq1a7UHQxWx
QpKLQJvZbK6LC9zp/paNmM2nvtTktc/Yq3rsRsoRNlHss/Gjx50eEfj086aE0POX1SLL4M8g0bAo
/QASjt6DslpST6VtgZxMwCiYNMVjQbEN0kkcrcm7oEhv+lgcKgOHLhn4J4j7dqyot/dxVnzuyIJL
0eFJBfkMhd6MKAmVvXEyJG0H3JhX6e8Lpd/commB32MMZfG5jleE6Nwath7fcomkVf5UOAjYb5+n
R5BtWYRlxlsIsBxFqmyR4VNpALcFHLUqm7ke8kd5acy3HsdFgN7kUy4xPZil5PG+iNTnIyUEX74o
dviYSClZqV2PaZJsntokPlmd0ms4qEorBmsnaH/C5ICN/Vpib55/WJQn5zqNMt72OnhcOMAKCCac
sxodca6SApQfha9oKRJ2ZxC7YBHd0bb2oASLqhvqHrgV5IHltMenqzkc5uNxFiydXXs5mdH1LuZi
kR/Vzf9XORdwURhPgHW7zBF9oRlQ+W7D8P+gbDd/on4YjiQA7ZYVML8Bd0ZYV0OCIwY7CFLlVEc3
ZGKBf9bAu9iLyR28ElS5+YnsghHkx+eoAfmCag10FNrSB1mgeLkcb2+oU0e9sY+OY70P1Q67hHh+
n5U/lKX/02s2n1aMcCIo8psl6ljUSRWijLym5k5ADiVd7+9Al9vPH7fIrJPNlq6OmYkt0rghBeii
/mzxHRDv5bHYID0HYXLA1QsNfPAuacSj9msgf6VI7aDDvwNFXlBvW5WN3ZN8a4j0gLR9TZpcPUlB
6Pe8t27uaHvkbp6mRslHEGiYyQ8UCIAuUfsuWK0AM9e/1cs9rAQCH8nIXcNmLZlk/xPG8pahy5kQ
ZVy+yO0DuKWsKu2zquB1p9ba5I9LUxIbyk68JIDhVIEsqkMsDTns3OP8ExdoqAnIdUZWR6mlAw/o
QPMRR99tIqo2ie/EeIkZMdJTwU2fSXC6UEuTIoZrGwtPohPl7NATHbiXvDgyV/AzadznITfY27H0
C76EvFtZHEkLHtUvQ2wbCT98ENOKEtKSZLFCTQruNe5Uo0M+bMYUGDj2ub5uNgDkByyfDzSCh+RD
WnYW/QnOXtq2vqv6P8aYcs3GqyOJVNAKIXL+nFXL3SC8ZMH6qnH776xXSHyXf91L+TH0ZubVKo+1
/BZaCN/KGPpMytXFgGBTv+NAHkcorflRQ6dCnyN3rnkaVCUpslvzQWNGTyeufrhfx5Bx55ySaPJN
7hbyv2d1MUFnLKGTOqS9qmMRZSVhnT2tx5vnfcVeV2SY0vwaeoe86bVsgZNdlDK/JXCpEo4YPzE+
9AVy8RD2LzyzM4pwPGWKjOyul+Cr9NJYbyeqek6leXSGeD5kg/MbhyEXX10EdbzoL4nam6q9uqC8
kAxMjH77z6OE6WhTz5r9K6wiC7f5t5htsvTntS6zGf/+f9yn+OEybudQajlG7z6K3s6lKgpZUpyb
6JSOVagXCnG23ZiAXXAge/1U46TNemxNkXQOjvmWs8k9VwzjgwJbSpTFCb3AyXgO5B8TaH4YoJOl
fLqbPygw+wsoG4xUndZ2Vj2gIPUfAScfvzEH54iOjHTWd9q4jRmT6lEfqSW0EYrGC7X7htqm0ERk
YTPYPi3M2FkQ4kaxn8/57gpAa0dWM3+d2gSw5ZWDuA4i5R1J3B8jrz9V09P8jyVXpU6DDLJ3mP/s
2WjznoYNsTvpDKfuMXdZpdk6WuEwxIIY0DBws/BIbZ0WWkTiyEWHsWfBuyvRH4XafsVnB0gbgV4R
vlx/a7xSwytE53ui3ZzjGkFL0cesRvGQM9UG9vyOjqqqBFf9NZAJAOP/VuXdpp75c/u0aL0ohEup
2ot+QWzeh4gnoXFfRibNaSjqg2vejtE5OHzr8JR+CNoC7aPd0k8sfJu458A53xNhtuz1bQcSYKrp
csnzIKiYTP5VTNOqMSQLSpVs3tB5halgdq2yLFH9vD3zFGj5Wy9fntxzSLlaOg6g8C7ne0UGB/uy
gtJAAz9NkVVHW+JphOP6ZGlN8BV0wGnCSNRSn3PFvLSiYocgj37dqC2CV59GUknddLwOl/EaNQtB
CKCuTybR+WJW5eBmOHHpgz5OG7eLVQRcrCOBsVVd53KdpAYkhEK3NBuEkjkb1DcMe4Jr05b09z2O
EddOtAGPfz+kieKkyYIWoLSu3qRFcNdCGBvAt4cm6DNiaQ7vXuig+2gcZeL8cTcrT5X4/4hSDH5z
9iti1osT070im9VIs0YbpdQZz1bVYbQCrAHyJkdYCPr1hSQYTbCoduTXfSU31IK1+8hhrBc8/2lv
5oZGA2V6cYgdreFC4RasjnkrsWGE1t3uanvz2f6vtBcXhceA8u0/bqXGylnOhmqm0b2kVyrhM7T8
0ITKnzcrBQXfgF3edTfrx34qD2/ZsdBdg8W9mRiC79YAQybEHIiUIgt1J6MFP3wbuBB6QcuIenJg
66i/jE2a0qdbA+Jo/tRRpzdA4ckqTqYvJohzEOxy78ykx54D6EFVrXnioXQfML2/nGuvtMPVA+fd
gqrOCQ+EXavbUNUYeV4T/r+DeekG2+zmkj8v5jqYwHdp/QBAh6deudArV1OKa3l+g8MIf8akMPjT
xIRFvNvgVYvmk3Pu/4CxTJ84pXNxZfUWJ+2k9hRMxCgPq05cA3dYshSoKOiWsP+zMBB51ZmtRrlO
89C0rxkaf9QsaPC8G6DYbvF03eycckRH82jM1/VuofLWUDOGRfVfzyiLj4t6Njtokgek410GB4n9
Qh8dVco/FH7H3MRJchwwJ83DUeOpGZQxmE5Gsar5jDshCnIeTALpQDe/naMFy97wgK9UDrdhg0ar
QwR0g+9VAbdviqhvVNllTfy5B9cUiXLGISmaoa0/Cyq2qrZQY8+fAe/IL2GRHs2d/x16SWqenEBq
4GBmBJJw0/GzQojlNIs4xsmmCELaZ8k00bc2PzUpAlLTiKHKbX/eXQwK+mVvKn/0d4tEtAH2zdtP
d0WgTHKyf+70bcC9qgZMGJ7LjKaCEY8/BkALEyKO76tE/q1iNiIYroRAZ23Vft01CxOkcfJSaubk
TpPcPy4bByrqFDVgx2yjnsJ7rpQYSPz6H6AfGmKbllaeDz2ycfTtM3o7N0zSWv4pNeI8K23N+ezQ
5QvyjTXz0utDQXN85u5WFHp8djYApFIdyl/ya3wsiHE0rGgsGGcTqSmP3adnuGLRzrSDMzB+MynU
wzUR9uEHuuE8d0B8T8Nm3Rwz9tWj6PVaCSAtnAQySYvGEL6enZ3MDQlwjVLjOOd5Z1Oq9pgWqmdl
3VEvp6Olo57nKk8UVA6ptkxG891Ek51hwaKNosc90jW7x7FT+eytvcu+02LN349NUaBBydolSqpZ
yAvZDsyjr0MzVnwOoeXK/b1CJ8j1wknvFnvOmzJBHPJKBzlxf7M9uYCBHfXG2b1bN/ZBNw/dcytc
061G05ZdpCRH7Xy6N82zzJnHXSfV1qWCc6AMlMBBb9xrGX64nDRPJ8JmjoACrs4DBDXGKyqaDqoQ
SomP0PHf1Z1Fo6zIboOWOiwzxpIIC+3C/4f5Ja68QiKBAXju1cawpljlsITMBhxGsiaUz9DxvbTo
mrI4Xvm15+qizwywxoQtEU5YJPlXfPxv76fzJyIbYxq7Ze9hlZlbWUaPO1ioeTGNG4yKG9Q/jZTE
u/LinZ6Vb/hfBXmp8J+XBwtmP1kdqFRsHmkfzsQ1isGz+JzjmUwdGeDuYw5kMqlnr1EdE+jOpigF
/jUmgcasSwIMwNHj6e0rRz7vw20SkwgfGMbBgzHsAFWsH7YJ4RFStL0q+4m7ZqpwkUvX/D13UdfU
pjtn32mYqpFzIewIQuV0tb90kZS5COz4YzzD+udQkn+dFKu9TxCqbjHUPFYUGemCv47JNFfmdvXs
mJvYrdUdHEKizY/+pJ3mgJlMnZap3lveitNr4oKpijfqezgfGuTS9O+6Qt03rCVK3yAPO8Wfk8ph
5ija2kheq81qWuduoQnjq1B6doBcJ1C+pJj1vkMRWd6hb/QrUqnks8fOU+CZjtETg1LR6DrU/pDd
r79VOOyzzYQiJ7DM9zaF926Wo6PJ+eG0+7NQ7X5dWp/xpefGqtE11xhRZRV17sri/KHn4zo+lDs9
yX4eXm/jMCp75//M7x2uyXjgUu8JvzQVUXDM6Rx8ZAskD3iUu41uMTYPQB0FqU2qhttmtjMdJDRy
POKxkJY1edqyoOQyJkjhAEGA4qAVH/rvIetSN/+NN80IP7sHDxdZKFvN15IeymHr7RSRU7n427Y8
3NOQkT0/R+yYEgFRGqStqwdaFdFlBgPJ7NFYcwK/K++qllJAMkHIoZ3KOcJLWsQ5GWvFnPOHAkLm
NO7ZLXTHQYsuWoefWjNLR9ph0+5A8HvmlA5VVvJKAtR+ssSOYKUnqv+1auW9/BZbGP+QudtSil9N
2AI/CxMXrnbEtbx4eBthb70GHyzJYzmqzw/6eQhJLkCPNvSsnNPrJiGGxAjq4UMjd/QTmiPARn+w
hmmW27tGl1qNNDaQmGn7g/97VUhnjqB5osPxZ1llgaEBfTStLrdHqsW43fLI42GyzHdy7crYcLYK
Eer7vQCJP8YMplA60m6i3NfPuUlCb2wuM0cjgBfaWtl0So8+QQu2ZWqHuXBLWXpqZsdcvctLF+vM
Leu3aX0N/95t2TpCxByCZTn9wu9RtBMfkDXjWgoab8EFbqRUB6BbTRHLWoNKfbN7Uz+epyIGSeSW
9uIbu5zvCA6GeGsoYy/35Sfg30nUYYM0PrTn69VRfO8QyRGV3Ji9/A/pt7oWgr1KxZFYfrX/nCZu
+ZBT/vhjlbscUpVqCN2rW7LLUTO4DaJh8ER7PIcV22f/kLeHZWdaH19szNR9wm0j6Fy/ezHICSGh
ACMVVqURfq9fG/RiiBZgaXL7M5v3EhMZ4O5dDP/08YIuyejJkl+ne6D+GiC+r9oRwoh1yGH+tHw7
lE0+fj6UM0gy4UkY1/q16F3Q56y4Ke+NdsEgIeTDQnEeIjrmXMlvDF9ijWGDuMpSRFTl33QRjcBE
xh3jh0aIztiU5YahYS9G7HJ+vNYRWmbpJ1B6Z1jlW/+jaq6zU043xSgv+kA10Tz09/WuZI2MzF+8
KYXzxWvi8dvVfg2SgtjvlLKpJ9j9423P7fxN0anM7SfthhGD4lpE3we5QZJk4puf67bgJtZaTnPV
WcfBZVm8gup1hUarpXsFhRGZtzYmhS/+KNicN8wx8e6cSOHuQZZpNnJuDCi1Cw7I7ZhhvP8xvZF5
H34UEVoosZrNXl7VJw6WJMOJg2v52YkBG5g9CorXFojLGVJcUD+QZC+eZeLZyBOMVyAVBE/LTVjq
ONM+4DRVKlWktsmzWQ4gvGOugBkCdKIhfKSQmy+SSXgjMFpdubKgb6Frflf0QCRFMBmk29NrK4XJ
nRkQ2OUILlkPG9C/qt9+7O0pW6m+LvRJNlT4T5grO6GS9gLsVfYOkSqFt5Wz59hjk1I6w9lcEEgV
r+YkcMK1TY00LObTbedI/9yQlZEt9sApdHFAXErL1rzNd6pDsWPmYZmkxKrW1y0DnVMxgpAZpyzB
tE/4N8nfgNIow0d8h6BLFatrxz9c31ZcDQfXs7JEFAloi0+NFKcM4/TG7fDyajH+Be6PVbBjE+C8
yKl4psCqGTUDDIb7hNMN2I1TuH+vNTUDZrLDf0BNFKRaJvKkAMcdsqJlOHbgNk0D2KFtDc09p+Yl
Zj4BZoJMgUEnMCwKiWql9pPH7+E+VLA9+wC8DAtw2W3eCSSKN6yyzX7aSKOYY4CNAA+UtpVz1gRI
GoGa0zb5gdG5l+mONc9xx9NM21IaZ36Gz4OxnqfZLtfPtKkW20QE1lNw9LzRSusHcMBSRhR5ZVql
W1bY2JnSojwPKJmWQf8i3j7/4oL0Ngsx32VSPUeK6Pc5nGnfeJTEPAPvyD//5BJ6f3k4fBsRZdbv
u3Si0QlFeXVnJMFYGT0TiC3/17y/xX0UOXksJUk2QvQLY02MRqgpYQhxipACaqGg9arb2J6ygFF7
h7VUK4fhZkVmvk59Mr7mF5oxaTZtXW8eoXDyw8uD3l5eQZnIZWG2Oze9vg1k6M4NKDVV2WheT3lD
8G+AG6+hAuL3JU8Qf89RGguOQy9KdfHgSi6ch8ZYsu8IT3LUlvtQWSOW1YJJ8neiy/JpjYduXgeX
ip3ETKLPhhWiYLBYFl2DEMH5CHUJDTVkk50xnla7C7vvsxztj2Ct0Y8AsRnEl9CZOddFgZEs9bQX
VOVKTyI9a8CLPvpg5fQF1ptF/nH2MZzN71hejRGXtiDu0ds6PU7nN3RYfyJsggQ1oGiNcMvWWEug
7gAbSfdNoenLew5R/EsczcpEtGQIeQB++yXIx6LZXYQgayQJDQiEbFdASLTQ7366mHwpK+PePdXR
o7JjoTYazQRPHyAuMVqU2Z6/8PRm1SKVhKTYxeE3VTHcDI94luWyGkycECRbSKp1h4MZXkSWtlTq
NhOP+GrzoCkAr2tVGhvBW2o5uY16n+1mD/pzyaMme3HI8m40p8b5WnKPaEZtRW9X066ZJyRqmSJE
Ansa1p+FMX1C5fRXMfhQl3snx307fefNVOvnDel044KajdxD6BIkoba4vJkJ1la9arjNjOZy83Qg
Q3tQ7OSf8Lkzsa89kJKsa5Z8ICAp4lZps6aopC2pg37tAkGSLB9cbGFx6DyB4RSvhbyfryMt8T+s
sXQa/N2WvH8e8b4CpXmaEhODdiaeGMLE2svYS/ZeM5wjsl+tF8IuzuKWV/LY5d9dCPMUXODq/a1z
TpJG+xVuvFdoxTIrA6/Dr+1QwMCqkknI5gWDgKHlBfLHujBauNhuc7m5YGEpUq2AQ94ZQ3jmAEhf
H6KD4T6KnbOE9QRe3PFihz/XVxBp+Lzu7Bi+vSK4l5ymdHj9IAv6NgwrLAam6T1wOzJjijMtSjiu
kqgVpg8DIG5R05LKpK5oIDN9lk9XVROy8gp4SrHihImYbRH8KIxrnJvpSMV+I3RAN7rzVVx3bhcB
ZU1ECJ2HCH3tata/E2t3eCOcCf/A9IAVN0cleo2vPEKLf70jOKi0TkyitIUCgTfu3SiuLjC7hIer
viXqvt0ThHoerdfx9synyIb1oDMXiiNwTL0QgeE0sud6wdkWSfegYQtPCTKQlGgL2daPH454OtjW
r/brOGDRamJrABPajf3Aw1dUuWhsE2sKAEnEHh8lNoxMvalC2TgaN/06XFh9d+4UotHOs89d9K3v
vvG1O8BmV2IDmCFfp4C6hjktsAOjebqaccuKhGqfkj15eTsLNeP+2p/3NPMMEO5gVZ0PC5md7CTZ
aiWRP4uiDyEB5t64tV2KvujpWI4+Km7w0sPzbuIoskESUbzPTIJ8zDkZbWnFfg5MvHHApq9iqB1C
r+p8ngX5gTFy5AwgMYPs/FmTAxQtNBIU9XbzTz1TrIjLYgBl42b3hRfrYrUn61kxeeTc9VY98dYv
CVq3QUJTqEdJ6S3F1CREz4DhDEGGqE2UjvCwxgehd4xi+SH+PgMZXWlSlViNANXH5IJpsj845u8+
L9XcuNW4lHJu/t+PjrAVOSeWgAYsGjJEfSmLngWTp7xiMCDqez20lJRmwkb4U4PGrM1MI3g0bqCZ
14ltrmCiaTtETgHHq72vaB41GLbf7Ou0J6ldciLOryZfykJOvAeqQha4YZDKLl6CHkqkmQF1PX8j
OHUxnq2j1z1cBkV/QMUHEj5x4m3+XxO4sFhG2xhjfrgJIXRubnz+MuQUv2nLuZXelpeK3UzoDV/t
FQrY3H6tLVIMRFZz+8yQS/wvPT8sWdTP+z0Cf0wXi0XjfIe98W1Xoda6IjN7Tujq4o0kT4/Ehr9i
XWXPzvsD3RuDORFAOemg0Cz7pncOVC2UjH2PidU6TXz8Zw7txZtYyz3D4e5p99PyDU+hARg2iK6G
z4wgw8fWU5Mh+u9KI9mcgozM4wB0VVWHEbLqAhqX2Q14iOCXjR97x6CdV0y8ts4Qzkw/WbG4gO1j
SuwWe1j1EFNOpY+1Z1qdrs/cpC3fF7fgIpP7BNP6wxJ/H01BS5ExEXVp2HXa60R7ldzASDraAhog
UjElde35iYAkSy2FFWHRZrWwuVliswZPbw3GujpzVso1QeNA5WbMZ4LL+voMUwb8CCnk8/DYSYo+
mKsow3SLM5MqQHwj8XDXVMLdwYn/LsDq0ocJD1i32F1YEzfjdmZ6Og9aIRo77TvOHdHIauyiMDRz
zt08cEpAtl5sJPpIz0f9uuh5U+glAwPn6SA3WcQpLRt8o+rIrltP3B8LXxf2dN+ZdxycxGAP1iiZ
gI6axTPsMSFWRxAExPn8p15HZVlbKDiNXF28XNq3WeGe7dHKXbwZjXi3sML/xY/l3aDEJqBI9ubS
pJ2Buh9g22LC+UDhG2GQBXRFr4wm/PgRckI80Pexwvsy/6QmxUrT3RaKMlUmHfaQvTnsPfWya/A7
Kyd+jrxVVpAHFUYNd0rX2gsPHvdXBS4Mi8pS4+V6kIEq2dhLbt4j4Z+9BnnZqUSFor9FWPLDoF1G
fZRtvbzjzkhJ425cWoiOSXO8FDSFigx6ShdvZg6jp9qMsIXKGV2exxvqIEunpM0vebHseBr+zlYp
OtZgS/dV28V3fs/CaunHfncWgl/lkcgA/1y5w85Pgc0jXPx2M4xMy/G8I1dvnEcpc6ZoMlqS43/g
eSep452EsqIagSEtcfruigfrQMo+f8CSnI04CD2REGL8t/SQyJC58I6yffnJmq3FHQM0g2Zo+ubp
TL68EpDaRBKC8a1Pu/FgerqwKyU4yBoRJRc7n1l3Ugc92+PYiUD/BZ774cg7ccJc0qbHRQhJGvR9
yRXLPNkPLUlhShgqVg9EleZC7XVM5NfK1PN5FMUqleyUO33XtYGP9zHMB5sOkcsx+Y0uS7b756/t
lzmx47dR43enN9pY3sPvI/yG9W9f7CMt8E662ynTGGErF8O+IoFa6HQS/FouUacnHuTZVrSl6mni
B0l/PJZjMSkykkgABG3FwhkiSnPSzcI0cHUHWDPjhkxSPWDz4XnvfyZNHekF51kllyrXdc1D4bPk
gxvuUtvXIK5J2nHgpJa3uY2lvHIZQY/4xK+1BLgpsYc/YOfCpU3jT6FITXOQBs1C5rXDb59ZM8aH
g93H1+0OBVfRAotZWMyAahanG/WhIkpWi3lT6qhRgFwU8m3g0BkdqrIB76mh+GwA8LuaNr6EUMmC
GPJY6iusAcgSekd/cMlRHQB0DiNTdjapNc1gJ6Y+ik1zh896wq9oFcurnFp9GiXVjK4iIwgVjqPY
naPavqXSLEBfo+DJUj5WIiJHnWaiKKfCIwX8svMQ5PqZDdcZ1xQhG1zdqgLUELeY6Wbe86rV1XoS
Q2Iv/0VBHmiZcE7gZF2JIRsX4n08n/oh/xbXWQXGzZTCC10utSBMQ1eAt44sN5pzch6xh+VjHlZv
cGi8zW9C6nSCVxwR66mPrukXiyKhQck+OIhZ4Eu0E3tV2qrA4c/u6YdGpc1xHSZCbLiX+rwmr6QU
lJxomchykGaqYF4P275UEskP8RrxJM6C8twBh9UrUWO0OB1mcM7nuMOx5EfS3wCLiRAzqLVTRmXz
PMwCkAwFQDN5YZIHUOSI4gXHldDiimv7mcy1Ane4aFdyj9Dn6UudagVx8ypc/nF7CBj1iDobDfOM
wbfxdAS6qna4/qP/6ivNU6L4ZdEEUhp9pZt/1gh8udcTeASMBWG+83rDH0HlAzSWozz87szF0K57
FMRj2aTOTQ1lbEeFPQjIO95awIdiLk15+0sbubcair2+L2vLsr96WztGi1un+jp8mls71Q8V/dGZ
/qLG3ZGEPCQd4eS2Virp+6bFbBJeqJ4efL5DT2mdz7m+/H/N3kUfWPFIPttALvHvD87W+byhx02J
c+Xvo+FK/OQtMtco4oa2F7dAo/q3cXBo4dBViX8G0kNXsoQroooesq3hSstXdXsEnHKsuceBTZ5f
kCcCZB+Y1ccrlnXzF5gZ2dQW9oFtOcYDX2AmoskOT8jBgwV60ui9jLrTOx/LIZaVb5/LVE3cKjRO
a1SwWUbFJcMnqJGRhS4fC9XPrAINqZc3dO9ognivH+ouMW39sN/Be/h4dJxN4gMMM6W4uOM++xdH
JAgaqOlxYBf/K1f/qPw/7MpFB9ZCZv9tY/bXVHgIUiNoVjAY4fDs4au0zo7hKr4NhydqE+iuUJGH
0VUogl0ZzTNkfVkg5jAYRl1E/lA957/mhCcBxTw0xbSL8FPeoO4yB3dqcDQdayTy207dVB5CF2Se
gk7YsHZylXyJvAaomMn8+D8EoeIL8bG4bYSV2x8DST96KJAzQnVrCifNunTqfJYG/0AddDpSXVSC
ru8KGjkDwDtAVAqdVUllA87xsZ36tDgpDyvpGUEyz97o+yCWQo4SCBYCjcpwZ2pIG4D4l6mGyESy
2MN363yZV8wDUI928DtbZv8IOCfKZh62tOALoH3wdGj+TvS+0evzxRVYBWeAaZ+CU6uzElmWAsjf
H1wPBz6cgdS9g5ztgitObUYOYVd/0Y8qeRx4mJ7wbvpDzeKE01YZ7f/BWOy3Q0Sm4+5p9Ffmqx+G
8gDsv6EpuvYKutEorQFs6ybsj0MJuqvM5BpeKv0rBuVBjp7RFSXidX8OeD1nTAbT6X8qUC9G+tci
oNT5q5B1fhOt9bn1RfoQVjO+bQklYk2W4FgK0K+9kqGePh++1ksx9955vXPmZBP2kEVySUWg0F2L
raLk2YLPnshTkqrXw2tUDstYd5HXTbTqXz7iDJAqDdUOkZEXE5BLqWjYdKmVdgfuMXD9R/smCS1i
i6uEQGE0GonbufGqMtlhPpEBaox6gXYZ2ynda8ASyO4uTsbEDRD6EZrh8Kh+bQSxUMSFufY/qNux
JlRzMMoJ9S/7v3BNG2YSNhsr74DnriIa0WAkqLkWmEaOkt4C0m/HqRipBp2fbQRU7xDRsgl6W4uW
nEVNFXigSQLywzmPp7CqluWXRuqOI6dC5flenprwRYi5RyO12vq9Wd2gh1usjM3oAvdJeRLkPeEx
/0JF9IdH/NXybGAtwiz+LBFZE5aR7AxTquEDM135rHPQTWzg5Q0NpYyLNBZRkd+R1iI8DKyFjZtL
CAzwm/EVsYRxeEO2rN7RqDOKeguh80v6sO2lzJFBki+RryaX+erPubdL6WpT/Xh66guatDqf6asZ
Fw8Eyfqd1w6yT+Klbipn4M4QWm7wBJuVn3gaDZyV11oPqiaMPehP9cT+hUkKb3o8LeyaDUpSM8wH
RRWLUHXcxJDry0C//7z0Kx6fg0wuQiSYGNsyMwkYXAIcmW1lSs5ChHq+n1QMaRK9MSNPjYqJwJ2w
G7lD7HHzCrAfGIuvoQycyN8EneW/xTM0HAnlEguGEsWgHI6cxhElQcm2vtRgpC46qDvDpBC1KXIJ
tZZ7Aw5CngpHDurfLnS8l9M5YVfc297Mv50rocH5tKxNrrpY+G2Fym3TphyZ+qJYR8Wqe0E6+6RN
UqQhhbWHCh2ZumeaXBApTAkArqs898vsPO7z+8Cxc0B2UQ6Ms8N26S+XlhFRYx3LOAzrQXH4JmuZ
+llZ5cgnyMqf539s2+x3x8CIhJykrsKePAzVr2ud1FRYrSytDVRIag5URalS/QouZLM9ZDzgLc46
LScarJ/HTP6RNgQQ4oRJHGjuOvIq7dWTN6rnoI9IVDciCIYv4U7my1OyUdGIpwE82h9Sq6xXy61l
R4uCa4Zd4ad6pdwxnxiW5gmom+aoa0FX9PMm9GPf2G4J+bFwHXW7F1YwQfXbYG9SPGXuUjqbjPiB
UBah+yj9+8QV5Vv5BlFgK+9DObiy47E5+/NUTteXxVdODmthNMQE+TuoMhaGBDA+ZNrUTow5MQ9E
k9QyynemCqRYUkP3nG8FYIbogthwJT0byrMwqT/j/3Oxmn2KzBOuFvehwN9cHw3z/+RbfbSOAe5H
pxB0Oo2hjFO0Ey4ZVdAyjY/0cZXr+DgQ9A7ENG6P3lJgaDLW1ccwVPFzDJMvZHyi0ewGm/O1J+EH
APsgaNjhIpFbNdiXgepR4eIzYwrdrJaxzAQ+qtRIMqvf/nJdtKgMkLfFo6wIsk5gdwDaDI8ED5VN
DbvWFR+73Hu8eZTbcVzakQGSvzst42S5K+wqF/YP/JUazDBwbGgOsw769OiVskhZxh1dCc5P56wC
GTnwGUP32pFea0El6kozn1C31VBwjhPzCBveKVyphDeF/pu0h2kzg+XZgRmgGtYuyfwO9176p32t
/MX2FYMVgGgzGsqbmZzU/Ame40v30QRuYlbcSqAbXaGQNYhnk5ddXar8mZJJNevtLKW09CFDst6n
+3qZACNg2ZO5TyU3XgvQC9NhUs2nasphfENTx2eYma3wvH1CeQq/GD2sQH8mUdpbYXRjVFY7Y1gr
TEZafb/3o/HsQ1Neop6Zl0yN+AJvGQ8IYLutXjBPr0qmuLylxfXbwGnn1emK2LLUUkRMWkfQ5DBq
w1GYqpI+RMvrzSWoIcB3r4hxmExxOLEn6NltGbnlLXHaXPKFc0aS+e9r0jsYJMQn2dNbiwftLFEm
Kk2GG90zS5M/qzwE0KFvSuWopE0HHFejkypinnJExge+FKaIQduEhK842VtOdCnD+UFGROrZEO3b
4XC62qUwDU33nleMbblPvPJKrE25kLFg1JK50FmNCDKW5HPJgUjbmHJbRJpoF1/RFUtsUsZMYo13
qnwymdyewQ5NFKtF70D9rPXQX9Mm4xwv8Zgw0AkUmpFloHsxBUJRlWpr76NLc1u/YIDnxVDE420x
3rVKItopyxKHMhw4Xbz7dqkrooa8Lp+PotXC1N/xa4hCtMdPNseKfYkDtpQnUFpL79N/Gcd1+Axt
gH9ywPiK+aY1+s7GptNaHml0BJo5WjALVPdE+bIiGg1Pcq6OuCJLj5fXYyrRgfU9c1sSl7VtvZkF
2Kn/d9xsvpSkZvZs0163k0VBwAmT64A06d/3Weo86wt1o1vIPgsBeCKDd93/j45G9K5NlH5dY3lQ
Eg2HlQKo/9M9YKGYD3jGaNl8B74HdHV8RMaDYVOCo9hVMYzifHLKiOYwNwQ5srdOtMNrdwEjzVAL
19UflLwDUawUNZgXvN3T+heVy9Mw3FCpY+dRM485ZG8PRFvPv7lJFaXVeSjRmzFzY8cG+YbpAXHQ
Gof7ZnY8G+kS0fvX9nu6TJkUiXL2GIdIHT8YP8r/MZ1KOygsLMrcFOprU7AhNap1QVhWuYyawnJ3
FuI+Q+nEMN/snBtTUllY1W4jVxNCNbYrbjeL3j37MAyHqvGXDIpf03cTRXKgCsMZFzpUWHvLW6Oa
9sye65d1lp8xrNGtwozy5bKyPdSX54VyhRG3l43DV/O+35CduddKiIqcPtfIUMKDeZrxMPu4MUwe
/HbisDUnjajQAmET8s4W227kUri4UWb6/6cH4/8S58ktpEzQSakDZPv+LCY22A/s1Wk3WyMjMElZ
1+vkSUXpYvHhx0aNPBWadu1X2Ur2L7JVm5SFV2elLq64z6/kb9F7DlWfMjy7pSeAJZ7V2UiiwmdO
4rkzwN4SIMoNxr+dRCVhXfetKfq07T30w3NETXFQ568a31aIwKLgPQvH+Jrd9reYRNDDbggSexet
hB8rc2xp5/eUVo4FOJS058tI8TCiuE7aPKK26OrHq7WhzoriLoZo2hjatRWaP2xEpwdgubT2DKwP
MF+KZIIVmd4OI4CSsti9V/KdQ5jjwZvXXCOlR8ehITOAGptOuW2dGl7Fqt8A6DT1M5plCseLxWd8
8TOWQiF3X746DA84rg3HfYKT//9+M0UQQbuh00P5RBewfjfIxADwmSLXKWm8/FCgaCDFwb3V6ZoF
ZoAqeIdD6oM2F41X8jPkH/FNBJaDdeOsxtWgjSL4ec5HHa9R13rd1WEgr7TEhX0fk1J7vxNl/CXP
BeFPx0fJT/+Py9OJQAT9nHJfFVfoC6qBNRG7bsgqQdsKu8oPsBNp0aWnMAHnmqlgYiqJ17SGSTex
ZF2IdFxAAtjOMdDtrZz2r3ot9DJaQLZPLZlsTFqqM1HhHBpcyWbbMPGxCR4x69ymN+XHQn/dBWdI
5WTdNG2cwwo7CeEOZV4Io2ZIJ4hv86GK2MLMgwQNVYEHmxvH+A05Q/MKA7qn0/tav2wgSAtktfBm
ajm4dUKujRMWeUDL6G2fWqrRQq19dawBidgXdojNcyNvjkTJbxzWRLb7CMFA2F7jzjh4p/hyZbdd
ghfOTMHyoP9x/+YPT1RtNjRycoVVsLYtBqIsqwRVp1AF7aery0UaPEgnbJagu2G8JosGEikxaDSZ
z3Jq41SxciRxl4mfhNT493+shpm5T+Pj0+brwfB/l1XOyw9vpPVneHKCN0AvMXDTFqqMBvz4uAnw
qxPWurm3/JFlY5YtPpvjS83ZyOlwc/DfREXLGvSpdO9VjGZt5Uod8WlKQj1zjq/yW5xcly+jXUf6
5bdACFK/bh3wg9PdE8FjhPwy3JsTfa83d84qcFA6gQkAg9Lp9c2qav8SWdppjZLVPGLQmqo9njNb
Q9VkGhzB4uePwmNTopiFOsgrYnlcdvSk5PpPg4d3ImpOUpcYF3/tuB/rGpthL/LXU7t56geIByKj
r7RQBk0DMTJ9ouEhTNZz/aoeuffTYBJxb/ZljkY3m1rqHdCyVoNkgAvpD05uaR2QeXTTEewHH6+A
H8tCMAbhW1FUuc0iU3hH2KP6gR23JVvg7hD/3Ox6eP+EdE5lk7VMqOOYLyAHZTqeUnqNR0AAdJVt
LaRGqapnzEUyX5wvWP389guVxbXXuCNlKGLfFRQQWnYvgUPO6p0OTsuDIj3K3MJODbg9peoqiR4X
CmI/xTT/4TXXJsmEVETlJJ6TYdOReKUwtMVjhSJB9Cm7YwSLmtWFYQ8EaEwIqwQyQQnH0RpA+W+e
YZ+TuVjP6mUBCqs14+nRraMSeGmpLIDSjVtuHaPoeuFGx3U7PDWHQGj/P6Ls450SXOARPK5OAj1K
sB7ZKEtqUJ5O/9OjKum6jKE4cHRti2L4t1s1la6QiKq7QuHqaZWkTsCxxUbnEMgbmpOCc5RcWFdp
7Fy8yWmwNFlkgAt8R+RnMByhpwKEEOwQ7ZxaKvEeqZMFx/cCkpHRFTQp9BrhYfkl0cLmyi5LBVdP
bj+H4OgF/RM4iyj/T892UyzGYeRYzyXR+1luvq74tMo0DoEHNj59TY8N4G5mCfm1JitSrIhbi+kJ
GEKZmz+XQVplomunxw/nAoScVKkLpBJ6F9wMnQpuJoIQVirxRLG3Ouu8RM4Zg/TvJ3uogGyYt7ym
7gaGsDS2EVouuCyWzqtHYhPtk38yVU069GI5abUJtLfJUjXmzp4qL5O/xJhzncmxQFyTRBbC8pX9
p5+9ysPVCQkDKHrjbgvjosHpm9Kh/MH1PV7ysovjRfzkRrPbMOfJvL9jKMCYt6rZUelmOTdTGC5e
4eBNNQFAEXyjvBf2mO6iIzn8HwYKTXMyzdUw7NWkdqAHiNlZ9HyHx4k52UM08tBuNl/zU0wCZreZ
an5ligZIC6/SkjDBqhOaGZTM6ROBCtaxYx9mC5jCuQwdG6Zvd+mQf/bZqa43f9UvWWfRqUP6JaY6
/mKAJGaDM+eZzKFkUigKNimteFpcpHSuc7S8xLve4cY5pz4bcHc/Q/aCPh97JahtHTSyjpAF0N/y
Eqm3SKAyawWDsK6QCn+leYL2liGaWuxsWYAHAnq7HpdsebwEt/ipmQ0tCR50X6uct2gmR5j1xhmd
2hN6baZpRFF51ICVF3fskhYM95teHHsj0qGn3qAEv4+bW5I7YKJJ3Y09aCjjat7rBZJVD+NH3mh/
tfkzdHjA3E7gqZF6+11c+vZS3WurobOdYK+XlXQDYg6lEGpO3twUjqNj6PdN0GxwYBbfoZ7OJnZ0
OTy61GpUrowHBdbJ4ojKKHlYyqL+P9RJhr46wHVWojHxUnmgPN64KrxoD729AU0slBGpOk6DHvrC
1Ukugv24j2UWxc2g2dXTAsmz0D5Usbm81+PUg+UIBfp0nmli/jLkt9rSud9kpCtvbGuJZ84GMlG2
fP7o8moEVVILoT+9nbwPhH53D3/48ubi9F/ksuUEKnP9XtIg5XV3k52w8MIvuRnbqODJ8tnG59aU
gqRrpvXPix89SdfD72Xaqd7lMKrMvDe5EuQqGSF8Imvwka8DEWOgD2CEVnqv+Pzqsv8GWXBdNbyC
bBnNq5FYiXctUvDfYrSSig3dSnl/dqDFyqjuM4MfDWicg03hr8j82+vT7uIpzb/K/CDmkDGNTYI5
netXlmpNaIUMpQT3HpPOEBuZ/+E21FL4iViwqVLpoANUpTbZtENlFnGxm70DKriMS6f4agoN7VLS
e2hwpbgS5v6FR03l3aqQnm9TR9goksawyPttxMq6+25d86cuctNGAltGHpwQmkBYK809KfOr0+nz
WRWTuecDZQtaOyi8c2cKG5cmDTwwN8KL998YCdoCrT5e38QQ/S8BbveSY8+n200etHzFF+exgmis
bVUwG3d6Uw1XRu0ozTCGC/dznpJh9uA4BZyF7Ps2lTL/6+4Iq6/q73618G3DQdjWYIDXMIkQrEyI
mAhum9InUAYIk8yl5/OO5ihru5uT54SzXb9crjoiipaxHGNGXi9WnGVO29tvWEaiahCrrMCZBTdk
Ks/hWpCbSmXArPNlSw6jeADqa/gFeOrszui7eNb0l00Ws/AXCfTWWqJgdlX4jybYQRwBZKGZA9vd
I65HvKx26964m/WzDVz3rEOk72a99cTJKd2qtKI2u0GVsk4XsG4snKa70/yolshIFstOREO1quXd
FSTRt1XUxnemHoSHvwFwuHtBJJUOJjhk6VBOR23M1lxqeA5P+Dk5mmfsw1o8z01TRHRyedxd3ioy
g2FCLfGXAZnYI38yBstyyQ4YIOs0usGEWj+j3pKg7t7kKLROPUaQT1DUXZ+qG3H+pTukCaL2uwPA
zWh/OLqxEvQMdeiomaEcakmJYWIFf1Otqx2vZaeF0waZ24J35H0lgq11w3xbwPxA4IT2lsTQ4o1/
cwHUyOhrlW3GVJtAtceTM985kRzFkc+O+jmBt7Hac9b3uEieCJkLySq5FA8RGNHAtMYZuKPhNi7J
0B8oz2EwDw1wG5gdEgNCcaJ9ovrRwPUcROgtB9tZN2LOV5Oc2SXsdyN4fI6Z4JhgjiflBqPJ2GTM
PyyJhiAYYNW61lEsq72gVHxJOe+6ZZ3zUHThTnzwE+Oxv+5HKW+LOZn/LvbnsuQnJgA2SdmtyrQc
4q1mQz6RTmadgO959lgn52n7avbvu9lL005YXKeY7TZgrA30k6N+A8FFkrRbPYfniuYned0bVbvu
Jt+G3epSr7A///txQckhdC6djIGVTQ/p4M2OAjTpy2UySZqFlpX06fsC0aE9LEAPLQKrKHhCWQg/
QXADawvUVbY5Zb5a5vjbmS2R0JTCBNgJAFvgSeeADmaY15VsM157XlSsyBuDoucOxH5nXES2hZIo
is70RKL7XDHcQbfyCGENUklpzDPM97kRItG1tYsp0AnZMtvJRSegbXZjCA/Bf+BePpJ9/NnvKfnf
ubdrdyX3pmuct9uyPhz0qk7U+ZrL1z1+suuoXIOigQOUIOy6IYgKGzHAGqfMXjyT9TFkZpj6080B
OoTeni814G6gKdbJMKlBputsux/AaceSHvar6DHj5Wi+rBdXq5d7LQ1RP0WV3TrnqHBnqzgM7KEy
8i0Fi3ZEw0xDmiNjGMKaJSo5y5shMIMrLH9oE7FbEvJPn5YRUeWROfo7LLuJMGIveqkhHurLYpdQ
eAqSViqKrXo1wpv0YHDXFWCXyEA/mDI4d6nOdHf8n/ZBUvAJz1MKmmYOUzJdt75Am1BTJ83nLrBQ
+lQH/Xd6oNlI0yfEEOq8LziT9puoCgCFrPg7jypOkVC0JBOdPiEc185gghGC8rq4K1gc0+H2pgoy
/oYI3g9fi5tdfpP+gcAquR8H8SfJKgEO4vtyp42Z/GlKF8DpWdoEop61GaczfGv0AU4x3mvVCGCb
UBpmAqnbb2d4OkOkupNjp5MH3ZFSYtdXvw/Jq8JmiLTiYa8XloAGsb7fhc8fuqZUq3RhnZcQrwoI
U2tIRN1UCe2UhT9V25dQScQDafn5LJxULIyb1u/w1+DTHVPcx9i5XhvlkTRfs7BzFQYLTGK/JAM6
qf7wqbCOYdbRqAgNialeeGvZ0S9iNSYMae9Dn+NKESidclrsweLDecGcExoLNxBl/yRofs6p1Vbv
9MvnpN+MSPIu3VroqwIrKv50aI16x8N6ptQXQGbH3SqFreDNgCyfC1glrVyAYua52J7YkjMdiERd
WUyn30ahcRfuRtY3VDjqUjylPb1w/MfVkDAr52mjcBGoorQMCzdprgUdFaeTBzNrC7UOWtbve4Xh
JhYya2A4rA+zOQGVMDpQrVKZFfK7A4VcKu4CR+8OaYiCcz3dkyQ9w/Rd+ulKlEvdPQX757s/cDmV
BJY2SMPTu7urY0qCTaDpDVB9P/8R1/IuiiBkuAHWRh8zGxol1Fdqxbblm4OEMiufAVbDBEAhomv4
UTPVIvmsXY+rXe3wBz8ykKyUPiEXSAAPUfweD4cnJ+8VMH1cO8UdLvCH4CNE8FkOPNoC8HPP2soS
osfD0Xf/6UsGITm4UBvvn9tEn+L9FB8smsrdx4c9VirjNhQca0jqVkVkOU0wQ8bK3JsSQ3UaZl+z
ed9ko7X85FNzMFQl3Qghvz+InLx3sjgx/VKlgLql8M/IyxuRCAyPkg93Gge5yiCwAIoXVhWnrnXv
K7HGo/nlJVyvFZY8zbffplgSLgG91lRJeS3gSUR7xrOXpi6lziaNl1eWZFJhaeflyoL1S+B9IyfL
cXHMdTykn/OsvUpkJddlRModPPIIDBSIm4PqJ8JBBaeb+zFjD8Qgjd3t/J3x1+ZQl+DUMEaV07Su
M/3daj+rwLAFO0nCJBV0yImMEL6VHNHfoCdJesBtx6CFJVflk4/MivMMKz5VydSWcZ8807TlvVDa
J0Uu2Yn7HQ5iPf1Zc+nhKDmnKSLxDfbV1u4PbONoiyY1m2j5Fbg36NJ52J37vlGFP7uKPfsuUg3j
mju4O5vjB/YsZYr4xwO+Q18Id1lRcx/hqokTwadViCeSJ1s/NENS2AZXexxJqCnvexsrpIqaGzrZ
LKsT9BqUXz8SP/F6sj6N9xqrumLxO40agKeyqP/jzN7qG2wm1O1GzW9D1cLipG9YEk2mzgjWVNf/
+gXV8VH5dN04vvk/bYX4B8xS+xo+tKu4pbQtNzwCHqmMpxpArJAOjMMlHt5fStisjWUvE5muZGuT
Hy+DVpPLrrF37XqEYb7L9YXBS7dN12EHp04KmU5FXYbmYcLgxK7VDK4IMqeWmIZMAr85sPiWrpV/
vKhXvlj3jfEwE0fDu7GKaD8wR5Owfy4xJYMmv43HdrMwcOJ9urJZnO+VWI8mQzRuh6NzIhh3wXZx
Y5E7d2rqcIwvj6DWL3ufstZTDJHhYerkNVAYIsQ/CUtajFDx8K1ORGPILY8wBRxR7P+8e0s3swW9
KUyl5FeP7xAi9kot2NHtNp1tq8rcTeUFMj6C2h/QFFhMSPpzCMmB5XHOq+X/+lypUslmI2qS68yc
CkkpJ5fwpuc4FSBEjqVS3FmdwwXt0QkX7SE8Wtzv3TiF9Zn0OCXqG6SUoRxXElGdkCNQdyzMvrQg
5VuEg0qOCwAK5tRe/wlOdo86iUWRzf24AG7E3oazqOYn96ttrmu5I/h8fbG3brNt7Kk1E9XYAc7N
COH1XguQx1LWYRChz+wY7nF+Ur027UKJsK83snARbnGqBzedQ7y3k66kobYtJOxv051QRXONsQxq
7+8yQM9koNXLJ8UERAElzxk5PD1lPj84mlOcKU5RhKU7h8fo2jhnXJQT8Pgsc5RoV84IddOPmUp3
wIBF+ghmnX786IwxD6eg0D1HK+NFYMoRxL2lOQ6qtBRSjqbZsvtOIBPkdu4SwA07khk5cBd9CeIj
iQLgL1/GVTMasSZFOWvVDPYVb+Bj8bVAMS4OyLMILLYtXPVHg8fpkUbekDNMppU0hygdc2D10Wrj
YGlTTFw049l8A7EMkogmh5P+JdsY+sbrzvwT8ROesP3zbvEZ+poygoyuAn7u9JZIpAXmM51zXHmq
BCtufJj3HBQSNv28FgkAdmVl8B9XbZxrJY3DSlsei51BLX/rzFVYr0Vfp2044psTNSgMgmZdRhj6
kosjq2VfJ3mrukVv3QXltF/pDKSxH4gvuw4zM0gKh0fnOGLlMFfE4aOZ07O5ggTeZMnxBrxuRky5
Zs6JTt4gqMjEz5+QVgZp8uxbFyMLup780w59sXb1S9zjG4IzHVrHdMTT1nA+diXOKGqe7uf38XOv
+LzAMowaTfWxoxMMnYyXRciOFhq1nmsjO55LNqH03LOODebeIZIZmDsaaYluhqqwK2dWZm2+8pgh
BaZDpRUVnlRc2mNKqlSqN9leO3SeP5mViBi3ig7Nk2LVbQEFqE/jP3bQbtUJ7Q1+1Wtczvia/NKX
pbVzG+dH8sMVz1Rlj3NGYiL8V+QYD309+mLTkVxSDISTWvqFNdIHO4PrIGW5XO7xXDAhWVGzMf4T
4PZziO5bDG+UK5joXfH+/bJbIXeM6tgGLUdgwVqOuJHsGTjNML5xX1x8K5Pq//hmyTeO5H8KZlQG
b296R6Tx5fNumnNdSkxYqUB+hYIUqCXK/9t2/wjm8Cd4lqpynCNH6D1xDdUsLHMr9Ahx3Ay0OB8l
TfDBBM5Oy5w1rF5g7B3Gs888F8G35Q+bQ9rIuC39nQqZiCFxM1OS5xlF5eozehK4egMNTc62A54G
670bzhsP6DCWGXj6PEe7YIjM8DR96qkkVjp3NzZDQgFPkvPLvmjmh+QqJJ/L8bIeJxtcK+3X6p90
8xQN9hRb+mwSvf/YdMGUoVPrpvEo18Ta/4J0S05bhhTzSkq5DiLdws18rRGz0UJij97hDPyXDHyX
yeMC0rci+NYgBkFEaGmS4ZKC8YtADZ3byS+ES9+iLxTATwXKcJTT2QKi934Xf5y/IVCSoRR7a8B2
mhYFFzKDFiPcb5/TNDKQWkAegYYGNUDN6erLwQ8u+IjZAABGIsumDVp78cKpLxzH/aqD3lboQwSa
4e/L0q93fm0n5m6a8jY8zlPwcmvmv8n4hWt7u37/MfTmg6GOJ08haIGH0fn79Fx/FpDxOuZo3j1Z
k6y+h9B28Wt0IIXfHeqgULMyna0En3DHnVnXCyylfX3DUIVuc0HqoxvmIqH1RaCoT2F1yiWzkTIZ
/QIE16hXvNyOxfXJsUGD8bm5lQnRzuOtoP2n9dT566PHFTPf+/Ge304xl3+op2BJcTtfDEk2rSqy
8LszjOOXZBuHuehuJyVPmJofbd1uW73+QCdScI4bCpoR0aBV2vdbfKr73W8p/qIrpwHgsEVpyxXX
13+wBjenZthhwFmS3T95nTs5Ak6ks+9HZJrcm8vmlWh2QWUDx6u/HVzW212CAMP5pRDWc+j152bb
K3lcUAGlUHB+TPSrpdl8Tg11sjeXrdsMof42x9oU2sNkwhlPx/EpulD+yTFOeADT1Z7I/Yoi+H5J
y7ob1o62HWsLnqmpGrKGWwnTXqzrzOsvMSef1G5rQ2/mrn4bVlEP59viXTR2XPuxXaapdbmW+/V2
ixd/eHmyjfd09R840C9l77zMisegy/dKszKCsUKK33ZWGB+usvfa+3DhgqSW5xnmfuFiJPIdH0d5
Ut7M5CoFrwhnnF9+j4L3LL7hugsBtiDo9cAwKv70ZeVJUlHcGY/C5DFRFbsL8wqDRabpfzMGB1T0
i9w37unLkqjjLFYQjR/9FFTkoS8qIUGZPw8fjrKCGQztn7iuw8yh/Wgt2Cxy/5RTvIz59vfE8VV/
gIuYrn2xwecThRMBWUAySkhGoBz6IbK8Tja6YUYiih4vwLvU8MJO/olqauu9543z3yT7n2DZXY/1
4nAHyGdxfvYwiPMChdRVTkPGCtlDiuRxTL+8gq4aK8nO8UaPNUV4B3ad5Q0aCW/G4IuumcwRTiIN
3ZIzMdFbGYSTAQUKPTqMlTOEqQZ/+D9gxK7USjwP5I6duJjjhbolcZ9Zf9zm3hfWdjwZAX9NQF0T
SLsXU+yHFsWbIGOdcky5kmvNiUUDfSqDNYRfsluJeRwFX5SO2nMRKzI5yN2+8RFZOEbfSd1HBwXE
1/fw+ghfem7POoJ7Yss8BDpRpdgaJAQU3Y5sBI3vxak7EpB9NByDZ7IVkJYHIAGz6VIVU4qriYz2
EhWcYWKzv0jMXrFGTbM2uFGBGpl8lJ2xXgPyTr9LyQuxFVQWlkLhpUzFYVIa9+fmkurhErP+eQfL
mbmjKsw+phnwGr4L4f99IANj8RG8oKlmtLXQhfWSgatcZRhzRNme/dUIWiPBAUZ3HUWjzD0VBhm9
Rv2DQMd5lltzA2upcXztbdmxmvYgsF9HsHqa+u3ETWwj4b2grVVLd1SM8Pl4MBX594drct5Qy8O7
VDKQzzo0LSXJvFXPB3m/WWRoHnrnuJilwOSXOlidKvffR795214PunJUIewuQV1dZOlmO8UVcB0n
ChFO2163a7q+SQxchuvU1rL7g/6ruFqz3Ff4oYBHOJpCA6jeixVnsUscdsYocv37tE5oHmaFhSzy
GHoWv13m91UCYQqoViZ6jkIJLebgMdqvYrR5Ph5oCXVt9xeqB856QtLLLkXwx0UK7PDEvndbq+ps
LAqAgEcKmpuXQEPX3egPWxkpMNgK6fH0jh53Y3i5j1nPvSxdf9kL4PHVe0eHqafU5hZRKPnfL8BD
3yHI9aCrV7JU1rOI0ClOn3CS1gWGMv9WBJOcGnn6WmdC8nBg/DZbtNyRNCN57T/8jFe9U4eNCc8p
h4iSO0IVKpMyruhJ1GPlgxJTseRep2B1f6JGGtnF8HRO30cuYOYx8WUVv+9rEidkQIVFFrLWr2sp
LzN5MPO0UAJUHv14WZ8vYb5bwA6fTRrF5nW3u4AhbLsIyYlXugMLX69p4CdTDq2t7aU2EvugEice
svD1cEKoVf4iehYu8ubPaYdwK+oZpbGa39rLVOP+7O43Yj3yNU0hkW9Vn6EhIEkfh/I9nQ4rUXol
v+DGyytCpF8+F+oTSiCSyE7tOTGFgeOjATZgojfYO9mC/Ot8ofmImMedmlIFYK4Y5FkB9gMDKUux
6He77/XPHI90lLI9bDa/T7O74J3xJjxgHzqfUqQRLI4pIdlmiMNMbbx8ospleUkp0oYs89lmybFu
862+ARSq+LSqUTuUOh4JLykRoVK5NKeq8330XNlzDvdftfe3/39HxuDRPJ2RVWpTztydkXprM2Qi
KodCQEXl8/0ekoWwfcpLyplJMkCvP6MUrxvdfTNNVNREzdMsBRFwaOLgtjkSrojCjYw2DrmUReHC
Mmhcdnk5n7p/Pmr691S/ftUFQXS1NHh+eOJ/TCull6WsmPwLHGGh2NdlHxDi0mjFjpuumIRSyVby
qpr9bvXhgPgkv9njwJqZvLTuLRpvl3yMjTkAthiSbv9NRjiUdjK21pllvqJdUs2Yvk+ZLAltHqNf
acMbWmtXs1kuAunsu9Cii14GrBGiw+0thsn+OFCUnLwf0bWGy1oDeyCs7vaPW2FxcwbOpX+Wx9oB
nHWLmaAM3l77XisH0FDyf3w/KiihMD1Pzlc8jTz6tcWh8QJ6Bgdrr+z+164cNGnHjnlyoFvMvAxE
Xk2WZqJjJIib8/rWaIemD7GmUHxky/FuxlRuZwUgeLDhUmXA6Z0iaoJKJsyCCVHqjQV7bChwWhwQ
UF8ZYZ8MXXpPqs5ApZKNEp1omgCfKV87Pswav3iUsVqMIWNma4eJzg/XhPondVo/Rrezs2MNgv7j
PvWYDxTjstoeN6XX01uc85L7pDsGJtHtPWiil6n/8sQCKYFsOWB8SF0A4f5+f8OQvmpOHE5uHFSt
vq4geZw75QwwShGF69iGw1NVoBLOc7hD1hrBhkukiHoAGV3a7k/APPoUV+qLpqXG1KpjLCCvpsnS
jXV4u5DOHXQGSIc4uoq16hxOP3mQLMzOaC17Uq8A4GD77QXt5hO4In2Ezbl+y0YzCHj2GqD2pPGM
b57i+U4JrO7igAkquYNFte1SfAYl8/19TV9MN3anaMFYyggCTEOEy/6pEqEQrTE9uPyIqAlCQsOe
1QWTS4qtB1X+v0Q6eOmOFuWfzlaXcFDtNBsNSTbuBErQgQ5BgFI7GkwVUKx1rrMjv36CibgIs5Wb
gdp19YUUpOcLBI9NliA4D4OZ6XTaaY9KjUJbwZ5bDnPEjcDfXdQN83/BvTjs06a2qK0w9XuU1NJN
imQreG1gTMoEhhYBD8XVvnAGOSwTadANrqFPzDxBzKX5evufPraWxIpLy4ea6lN7seLutWfH5mxb
y3kqRGD9TZh7Bue1kL22cNAZ5VQd6y18qbs+Ujh/5jaCEHVpQL3MJByAwqP7sr3fdmmPqgYLlEAL
tz+LwTyCi9u/Fxmz1NvkbkY98MXPmxOSr+JOLG15R4JtCrV/Zg++3AE5OtL2C1I7Q4XgQ07bwI+7
pMI344SHTqABbl96fI+we2xZeqomFfxztwvcVJomVfrL4ZKc7pg9UGL8Pj22DgIwuseivdqpXaLk
7BEkJYG2CR7+Z6ZJ8PcTSM5+LWcJkccqnD4L7CXv0Tb7V1Z6IE3Lnc2YeA4+AMhBpS+F6PSbyWf3
4qN8YB4eGk/7QTgjtu1DjD/UNVG96nwBO59aAO1S1m71A2oeoPo8qQ832pqi8TBxuN9fWaNAFSks
MYjsjhS/FkPB7mMeZykoUmeVS2DCw1UaaWco5njwl/ahBXJIv4pGuxOIW+XqhW6uKPykK+mrUw+k
FToxP7m06mmi/VzRg/0H9QfzUWAnS44asMiCufjVq8+U7xXUlpfbwOLG+PNo5HosVdlB+Y9J+nUH
LHtWKEStCf3VcEfrBb37+f99Dv+hiAn6Ak/ri+NmCJiYOj3ZauYSMbVQ8zp3uT8HyHjPTr4/5o+Y
uzsfxG8BMR6IguxaMwj4fgnlqRaVbONoWvWt4xhlO9He+HfrLZ4Rs90V+XllurNoaUAA/3MZ7g56
Q2ezkM7seg4lWrySnUOfPJ+l7E2f4DfxQIc+je9CSMBq/AhacfkS+Mgi+51xRcn33lc4WFIARSRQ
AV6DONinj5DaA0+1B94tsZEkErmJP/u/rujYU5wayAvIA4ygfWXwepPc/sd7yCljFbuIWH8A1B6/
+POw5hqVMgHGHA5ukB48i8GJdXDNslucS3SGh80TSJ+BveBy9x9EON6LXdpKKP18Sx9yOPqqQhMY
kmlX1kymFeYAWMSfd3NoC5wun7CLWPTPnB/UQ+YD9uHRZJ0kjVgY00V2MW9UWkuBv/IePHY2i/bF
lrSieBk9dhTYsUKLMc5njiFLTOZYXpit5ZJHsrLSA9BcLTM6FpJ+97kaP7EpcaNCIT7Zcp3AVJti
UG2pQXJkWD94u7oj4AQAnSMWazeI14tRgZOXyp+An6uztkoftaQSBENDlr/Hxce7ZCSKt5nQ7ngZ
bHy2iLarYeq4HueV0HObu34/lE4KllnwankaOe14rBRviOrQAQ86zmlcSqpqM6ShsOfQE54OtrQV
HUMq1CaxAA3iXjbZrNdJBR+OPjIhrFensOGtwKijjpbq5ou+qWQaDNRKrPEJIHhtFl6UYFSujMcd
p2oRa3vOpxcTND+VhN70edSQK1yrqh7ko5NejAJskVkiTQfsQlMLCLYunV5rr641eT0c86MBYJvt
MYP70Bzi567a6zqgg0LgpmDEumMZoAHKEcTspX+ev9z4EWBuO9bGCcJ0OE2v2VLBHkgJcAWvqbX4
7EG18/WaA3zdK0OWYXuJmhvqNGDCCHaw5jJo+fQl29cqXh4ukAmKq+zCt6CSnvbNF+XHyg9qMiI2
YYMnFbAaSY0KUoZihHU2V//NsB/Y/OXdzakYqGymbfIPYNTUGHUITuwUnTOB6ISXS+pUGt3UHe44
2z5Qwxrt60FMN5dR+kHM/KlKH+jrnyqviJdMkV5grNu+S4c8cQo2ytW0I0lrPdmZvZ9obr9SgwMo
1FnI67paTtSfQxko47t+nEedvSY9m2H/mQp/WqWN4hP1Siox8Bw7T3Yn2iov/t78AEz848Iya8g7
4gACW6Rxm56Ob7HCQE5IV91Jtjg2N3RZeoQV3XbFgrBe2SU34FbKJMxcqkoSUU6fpAF0YSBuw+MQ
AAy55+o0V/y6SZ6h2osz3v+7MGcPGcZ9WdIugNgldqOyp4G5ltqFLqkXGNoVuDk+BhBmpEw/QOCu
vhudRnClwfv/cLlNdPGkNregOr9vzQUbR/UIuWeRmn3kdo+mtdeY/KPTYMGO3IR49qg0G64AmuAd
mnrZ92xeg1+/U5ED8AVY+FbVl+zgsSbhhTvFd4rBEBNFZn6fY7taX3bTi66VpUTteiu9WCKQ0VNn
5MQiiCYa0rZEzXbRg+xqLc4LkV43KgftXePH5vRq0LIrGPfDA9T6eEj8kzSRcYPrmYo5Pvq8xM6L
ruBlo8SqqqjoJ6w1N42iKQ/D96R+rE+nxbjnT/SrQWBqlkWw/Mm1oJgGXOUvWXNBsgj0MCSd4iMq
e+Usu0hI4wM2xGQB7/D9uW2h2CCLRnCVg2ab825vTI8Re22WEZB474vFAkkgfrc2KBwsFofwqk6q
VoypG/UHK+oE7+jbwloXWrPovrN9uRlQgZCXFr0BFH0DXNZJCYZ/Q4JWJ4qNAQ3i7Wm/D/MB53jf
mNDlP3rZ3hphAhDvgpeCSqKYHr/vSIFgsoufwLFsSGkwCvxLetZAbtqAXtseaiasUX1amlckVfZ5
SzzJI5Xpry62D77Ui/8OyH+6V8HKpQs8gbSvn+XLbRq5icEpOzZojujkMWRyoDuiPxRaVVBzIuzP
JBhUKSIRSOQaKrpaQj4Rx+iUR3UvakWXqS0hXvP0DR2Gexf0Ij74SaHrnNZLm0qK6eH4kWDOZkFt
l4cIqaRBUBBdOhyvtrAtGVYPNI5rSlP25sQ+Xiq3QsqXxycTwBakUQ/QsskJL8Ve6kgOtz+O0Ut3
rKgCUKGrkbAzkpiJgxHJADmJLu8qU0wcLlFpqsbEqXIxVJlbXUii6y8bUf7sWfsP6Q6PQqqcwNk8
UC1Sqouwb9+UmS+oWTuYGZuW6SGkvJnA63eMeDTppl16QnzXCdWkKwBPkOr+GLmEHDmLuSibimnW
zpS9ewytPpcLMQhnyuS0RggccwQT3kKhH526tpiwBTbQ3/w2xOI27oQMpYrE6TtKhlr8/XmpZuPj
O0EhZaS/O+cJOttE8ZptRB8AhqpW/7XgJ9wovzVDEQrxakCWQSuRJ8/nzg99BLoDz2PCfhAFKzaA
tlHgsDnk4k5F5Bm8yprDKJigPrI5e6VcdkjfXSy8MhdujGGhLbnvIXTlinSpJnNvkkRH3Fzf8OwY
P6mhgHStdx6evkwTc2cHUVk6oIQls5W3gVfyLIYlv5i359eWm5FxmzWbaiylk4s/kWhqmLSsG9Du
8hwoMQ1oGMD5onH3Z5VdB3zimeZ5cuTVvwEFLy3gSd5xWXTXgdEMWr/EpUbsK+Q46QDEmcUlpy8A
XQAGHFlAazeB7knxPHcDF7PEbNQj6U/p4dvrEXsNkRuUGcsS2vQHMLncMHo6O/xytVj543dhzT70
by94f5FDAhN501o1JhWaceMVHaOVfKFGKB4gRnf0pwTGzSAPp1nSHDrBtJgQzihXZBqB9+v7GOf4
n7TF3RMs54Tbk+7gGFimCsVd5xiAX+d5Y0nnQkNWEFv1Z63+i8jltRbMhW+BSe11nGDz9CmzEdxx
B8g4Bfbrem+qe/UNqgmtzvb8Ax9Rd8sFp0fqsFZPkzTWFi6ZbZ4MbJMkS+ip0+UQ2xEYsoOcKLic
Khkjy57RXYjrc/sI9eyDY4L2c7L626eu0udxl6BnulkidQocxnv9wUTeBJTmYPtObrE5W5dNl3zX
C/RsFtlItggoAtzc6eLU1BIudXZBx/wi3vnrHItYRF+4Sf9SDG4EZihv/MINmLEyk/iR3ysDtin4
XlI7JxEv+sjLGNG+YhT+e5udlizGJfiZk+sSaGy4GWnzyjCXeEAE1EvfJOVcJ5F32gtHGKsDjtmM
5hbC90X5OekTWRixZkX/qSaNJxWVkQpL6xU+ff7mUeWxdD1tMtDxLKY3Aj9IqgqtLhzd9ILN8LyD
OKgw9o1N73xXk1N7SGgzvkIh3nebStoAzdHeVGewp0hzNi7vLwNx270djtz3FvD+4khJxoKr0CQq
iyGGtjG7TZx/z9ka4AgF8iAk6ruEBOyovemcqaZlX8Vgb//DNI72Ue5rUsJj1hG7MOuBZEMm6Xpx
eFvjxbIdimcO3WsGiDPY4GcGi7pH1dSKA4W5dx38CHphtBOBAHOoWugJt4NTZShziI2WQ7f/45lA
RDK7ifTuWL+H0d3W6SLjLELEcL8hUIi+GXZQe8rnaJb1QRFdMHY5vTMpBwGAlMWfHtPc/3KzQnVe
RJeeup8JaiXzGMPDzzbKtGBP1Y0Vgq3zvPnw4HG6PRnuTxXLIi59GQNj/sVw8JE1M9v5rU4MsuQN
wvDopcLBjDyGv5u2Pp9kVILdnA1zufJr5LbiH6cN9xZu7Z5Y+PHbpzL12Cl3zCED+imG+nvFdB7L
78qp5YM8XtjsG/aTU3q62M3YeCW9rvgnrY1HaFoHCLP46RNGN8C7q6sfFCWy9ak9IMcBVIFdg1zI
En/BL6NmxYP314P8ddjaWU0MMadpJXpxnTA5xLYNkHvRw0/Z37OgI7mx8Dc9jsJKh/YhhVUAifoV
tRq3K6sWQje+0C5Q8i3gW0oDMqeIT2uS3Y5dXWRXMc3rCq/SDa7q4aZgFuqyWfBMd7q4eZkXRnLY
NA1dSYvFj8Lb6wTPCNqt4ZLiWhmkJd8enKqQqU50pBRpoNi3PojMYzFE/k5/3oHi8E9xBEEsbv5x
ihHusQTakfZJ03TthXeitRH5Kz/w0mrMDVYAVx+UwjVmj/ibJtkO8fR5j+g/D7T0uH5mGNReBWmG
a+Fchc/uZL/TdH+p1ARnA04LJ2CpuFsXeEqXjtJjci+ePZvY6DEI0JQlK30Iqo3LBOlByXoUqFGQ
5miBDtZ7P7/awH2RRzxsh3ddm8J5iRR6rBT5Hk+Ahc8tbHSsuFCWCKKs/h02YYJHJV8GLMcq+KCv
axAJO3kJTKcumYYZVF8rHTzJlw7KG/hSqIqgKMEmP3rSVGmMdzm7IGE4EKFtipgyFLuygB+I0S4J
Cp4jI5/LxA6IeuSCHFB2otpyo8aqutCe9MOu35aFDwdz7NHQYTt2R1CT6U0RmOc6qW9VkiVgsePo
UOTGtPBY3423qFnFXAeSFJgiMFa9XHlFR1SWVkY3BZai8SZLUuDKiwjH/yTOkxkoqw1+CtqZGU8q
vIyWmChQTS/ntckaJ3Pm0Je3cXA9XMJMqhsgjjQI23ISi1dTS6PUbQrWBF2t25Oq4CZeJViNvLkn
ZJvZwUPPANKg+iylW4zavUBXh7X+WqSbik4SGxfx6DYqQc7lkERZOJpQNlTk6MiphRxdQAMmNFdj
5DCO5cI6JxAgVOiMmwikLc5uPaGy1Ltr5DKapRxepav0B2as3pyuOIKuHMnEwA1lmW2+3qpKylUA
0741cgHlKkWeImrcAabnWoH0W812zkqY/Q6RzdehC3VH54d+kQEaoLoLM7yUGaeDB9P6sftqKV94
oVdMMPp7ZyVOSQG3e+DOp14I8FFMnMX5KoyjZ5QTZE2FoUo0OquLUvNTQhA8/5FWus1qlfISygaD
oYXzlVCg8DRMtuUy2JlEy3qVMN+5ABKENV6PBsoBpWJWQaGmBClstfh1y++NCAr52F277sfpJbAu
nDWaJXOmD1CylQ7DZs4CO5eu2JahUPvakjNsYVi8RqWaxo+GcSvJpco1hyE9vdSCYainnkaAChph
C4DvRun5HbHJ4s+EMYFqI2weJSiJtj+VDY7F3+M3o4942sG7i9cZXQ1rVYEm8KSuhqhQ0XQDZme1
thbTfzzOLAGGw4Ak49PhSvVS3gXEIDVCZiFYO/WqRUk0Wp4dx6FvUhY5AoK63+VPEJExMCtrypeT
8JCzqQtmW29mwS2wruOFujYGpZ2awddSOJAC5tNtqrmyvJhVKrPK2e209R8x6egmEoYQzpqhIzAS
8u5uBw8CjOrP3say7DttyOftqG18ML0xeKIwT1tYoZ6Za/D0GkH8iH27Uuunp5RN6j6hPXnhsE5h
TKFpqzLJqDwabpz1MxAff5fzk8E5Q1E8Ha8JhtIRPk0+1bVI5uL6KwpyDZRb5OyV+cdLm/sIiRyc
1EXj2yH1tHb/nBWjKKqNvsRyDY/xFha9wg9Dw2RAYN/v1mjDST6IjzeiuNj1d3T3g7HzVxIY7Erh
vA3GHeVRtL3R+TaxVAwJchoRRV8O1gFVKVrbVlCqR86ls8KHer4j3QkJi8Xu5g5AoIEoJnzPaoP4
qCZ+iC5f85hem6MaPR/IsSUGpus2raViXF0jhRxR+TrA1yLWDDEV5fhOk9wn3jA/0JJgGa+xxghE
QTtNDYjA2r9sVlmLTasZzbTU6czQwAHsodur9JsRG9tDBHFRBBbjb7yGi9cdw1pvT9h9gJiDpgV3
HIV1kg3f1GVYw+4eJ2GIwjqFbH/1Eo0zX5DFyqsQe90mpqemySW6dWcbITwljIPsTZ3+LN6N50A0
4IhBQOr/xNwh66eVFT8UkhCYG2pujkBZOzrHaQzMjP+Rw4tegXkpQzuqjIC3JijnuaZ4+ITeIzsF
aHJpcgIYVrB4yi5dDWZWUN1oYYpjgP1USa9Qweyr27SJv+iibiNdtMgrb+fJHn+bV2G+ysXvr3ar
kJ83fkfcRwwVbC6tMUx8dm01OGDw8P6c3JWicp6WpH/zLANvZZSLv9BS5pbe8ttJCcyhH3CvBUjl
qi00Lgd23L2lKLDKcDuQ+m/oT9OT3fKbTscLHAjJd58KvrgZfiCTV8Fjsd/qg/VzF0kfS4s35Rv6
esUm1GlkIIxXseGLZliTYFhJ5jvDmNZtDNg0cAIVWwY8HHnI2a3kFDG2CUMs79BWwrTzxcPrEisN
kkJC0RGaZw575Me/kMZ5+7TAnjtdIlrB1iwNlsmGmA/RZ1mvxlM1WOLjuHfULq0nKmfkEOUy/AwI
jqZv+ZBeNozadoMPgTxzYWyGKK9Z+WRBX9cUGkPDpbD2Cqca6sLm4FPY1ujko+NWg9seC12/0ir2
AivvZu66pBR4RN/NHApIsjkC17kQhmGS0oEPFH4KDqc3nk6IHzc2rI9yHMTa+47GTtgCzSrjgk0+
qCwrqcJsMgpJuLI7wV4subTlCQqrmQEdLglvm7TyMnD5OJewkTOEXB0gmjScHAbEQwz8eJLZ1qLY
j0MFnHcRUTZso/uvdri5MUs9ZH0iyTqgKfiwm9uSMaf8c9t/CUXW8kNU7EjJzcqr0PEmd7z3DmSY
PcF1geIwpY4Ttj7y7OlAtOMVGlUJgNoXDTpTZZIQXo74Dreo2BTPByRfkoWF6U+ZOQB2KhqUKeok
sHmfyjHibWl2IYZ1yUhjKaXFlbhpwMDA41O8jZeFW8DwXXA1n27GaF1Ey6y2thEscfY+hVqL/E37
AX6LQmhTICOOs4Mc67fzo1ZNaFACXEdqLBoX84PS/U1T9xpLA9gdMyOUAkOGjsjhOvR2wMTBPzS3
salmkki3m/do5FZ3nXmeftMAeUx6uCTTIZVqPt3T7XTO1H2SxN63/4VOJ0CtaFo9ni1OzkV65oj3
mxyhZw7RuqLm04bI3c5NlYrUnxW36m8gxSu7sk7QLVLCYgON6VuTEgoEeTCVVWiKweWb3lnKjDf9
BHXVylNi4NjgAcsprvnycpS+jOak+FfyHNl5sYz5I98HNQAn7ZS2Z15ODiKuuF0TomdJh33Uw4HE
bUktUbahMsQrTOI4U7789uInYDWQavjrds19mv2v2I4aI4NibINDrCGmhbp0M5vQftjX6Lw5NvqN
PnSriGmOcZ5oJPzPmxUPW0oyeQp18IrEDDGe8nScF+Nj8zciWLMYAJZLAaRZ2QT07xIsKwfPlt10
xXK0hJEY5/uEB87oLFi/4QMzDqlLxCvYs+1Z+TKmF2+Qd6B+lto2CQ6aqDq2GgXH/Q7VmI5UELbb
WT9TzI47F5Hnbwfn1YN0CX0GRhCBSxL5sftORRd5+BHtbEc1Lcy0D3AVqcM2cq+lcg/iPX2iwh9L
n7zMmbKFJn4Uvgw6AsdxEn43z7UgezbIXN7RgpU/UbqZliK6eWgyQbs3I+RL4JNG8OzfMP/xc5k6
Z9U86oIUXxcdsOczCc+fwG4TIGCeEm1WKqrB6U1FkDOydlAcWF9p/gaK26ddf1Er4JE52Fc1kl7D
I0DSe9TtCQ0aIsReAmskoDPAfGdZ9dEWlcTp3hFFz95AUTMvpDIEkAP6PSowF/QtRhIaIgE10uLx
/+BBphbTKGLPMIHoluiLXasCI8eDeGxE8A0eCNmJlXZO36Naweagr3toIqoZDH56zsDySxxCbM1+
Uwx4H0RDuKzsxaxfScG3qZIzScF0D0ZfwcD1BQK+GgiXLVnOQLEmG6ltJ30HMDHq/ID9Fd003Mj6
3EKVNshiYQ5KQBc4h/T3VUVdN1JFDk771iyhwXjt8rSKKaY2KnlYEd4FNN1ShXZdPAdZnCNRaD5x
qsPENf2gcTkgSr4ZRx1Wff84C0MfiTRjCBSypAUUIhO8PSH9cBDIDX0ALpn4KEftyzpFDqUoG7wG
PVeBVHiOl6y6WYITUsHAk/qYN4pJ66tTducjTIuDIG+1rUfRhV7mob+ovo8CvmmWX9rsDMx6T9Ym
/9wN8nxNJ/dtRx1qaNt2ODTIwFB2Zbz/rk4iRXY1TbbZqoxoaf6lJ6zeh5NNg06s/DcJPV0hd2yV
YhO8QcG8yg0M3viKEk9pMyv9HZLJKlO6g7XhtJTFFb7MwrmxrtrwKEJ/03eQu9SeIlGd1eOCTM1n
mdFyKCBnQPIrbBwgX3MnMrQriEOISGTrHdeZLCAD0WrYwyMuWJCHalq4VO09tn6HSPXPakXT7R4i
JPUrwNSOGJ7SFPEeSw2ia9a8JmqWPrXabT+IJdiu1+pHytP/MQVxnRnJTPlHSh63czcbIFWlz1Uz
1frHGr/aXPKlXpuxajRAFifJWwLl0crRothYu/vqBoHQ3Osz2arYGYZfiUJlJnGnqKCbJh1rcxpN
uPrt7ZAPYJDfQHTqDfM2LuzfS3Gxi4nNjugRhM7fqPm567mJmWHnH5YyV4HJH9CqXLSgBcbNoATK
0DZhMvH6yL5Mydsji/QPaylfXh1E1Miqhijeqz9eaw2z1u2EDBImbraf3dAecDwo3yRcnbMC1H1p
OnUOzyyINqlDah/qPIr/VnGGktkt2MvgeEd2qoUMmR4AMfrZjj9B2Nsj9sXFnVMYQEz7FwyTO74e
yKkvXlZ4O1wIDJaLOA1T0jMnxlh+btzPfQOP//bSiThwZNAbr8s5oxH7KM8RX/x/BQm3qO3YtuTB
U/V2i26RNmKOdITCN9+LUysbEFd7NrmeSMBivNw+yaMXflebLoAZIQCj6u8IIMfQxN4yBl8YbN7h
KLXcDO23Md8UbEY4wwDR7A1N00N9QN7QKpu7KsnwpEmFIr6vpjC0l+vSZtDY8BtXzegZ6bRhfmVr
HYoR3XFkOMd0Nf9l1qZYu8vR5VBT7ij9pTAVJ5Bk3usx3JDLejWiKvFjlLy+TSe5wExvcEuh9dZk
OAvPCOCOf9+cQYT6ODU/sU2lRc6zIdrjcEgskegcNXZ2lMfVOpEmfyMocANCBwNKtdpIgNP3GtLB
y/kcNYv6RKpFawx+MiA6Ighu53jHTda9W1V2KOR4on8C73q3y3HICCevSTfJGH2kgSis0ZY59aNO
55dKOL3T97gulQ5aXBrqI4dKrdUPA7wESDkJWpUahPE567sxItDY24HQorQn8vjk6ydxMAF8S981
C3GtsLDGse7Qm6RQULBacmeWrhV5m6BlV8Ia7f0YjRKdl2AapeIvNp6VHDJOS8+x24ocVl6nQDQY
UldjItb3NjiEQ/rMAZiDmVdokj1HhzgEbtGCkKx2QO1jNE+OjRpAfuDZ+evNeVE4EiITuS8HSfBd
KwRnRSKV58V5ZVzkMsLuUVTtYo4ahqKlEMAKaW4le+QWfTG0+F79UoF0W+NUnVITn5SMHbqPTXq5
FiInUeqhciGQLi+KB6gpXgYtaFXfmtwVDYihmPRNI5IGIrkwWe9QcmVvJNWbM/NamzGcY1EyyId1
5jDY/jr/R974O5h7Gtpw2RljDotzBLrVkM755/VUDePOhY72ibsIC65JZtj0/LTxZDazOY1B+mrc
YTrgJhzr0BIF8POzKjOWMAPtf3EajTIllbdcDOePds612qtn8yGAig4PH8d3/kPinPdAATZbldZ6
lH/d3CaT3s52DTnvmgO39ASO5P697igM92mzLUikqx91pTsxKfSo5Nk4Vu9SSLaMdYCe/vxlLQBi
MlPpg2Nez0fTDXEsX25YS6ojDj6AMkMQ7YKf0GqznK3n4OFemfAmk4ZmIHLmjEvzx3nhH0aWJ+DD
6vgUSIzgJbvrm9gAYf9wSKiQIffL93RzW0Lq6u0OI2a+aeUH3zEaBCB64DgrpjNiRLq2FY90h5xU
LGK1bGrInAn1f3VAefEUtJeiFLEl6D3V2wHkP9JqSSbN98cvlB2vyKYC7zaFKsRHGRNLlFhVVMvd
0X/67VpE1soFMJQTqHXwyI/GbFDe7EJNNqopBo5sFZFSUmWm6yrOTlhoRTgVdpbFN9bC07RhcmbL
neewJiwz0veApV2p6YeVTlPTvMPANPps2i3apt3Qsm+9kFZUU7RHBL9sgb6PXqtW39F7dO2GLckE
O2KdIK4noj0pEBHWh15Y9gclk6oFPmxBTzo51FFy2OjMBzslIbvxd/UVmw4wWlZeIUooPHLpznrv
KRhpBftWP0g3IxOK3sr4BywH8aQaBSWeNtGWM8qeCQBmmog8hStuwSAG7VeDxPtIcwJc13lft3ax
LFM9RSmzGrYQBS/eR9n6nRuw7d1BXUj6+yfHSiEi51eScXIHOn8TGffEWz8B+htOagcoJr+gXO7h
aIPubMulo7u2VwGaPaWVlqkVJQdG1TeWMzT0cfgjiym/XdcIxxcnpQqwRDc1zSdtyM3y1ycuej0g
ETddTv1vMZ6VkE9DSSX/ia6Hg/BAdq4FBGwvxNvRkqIDHQ7peTtCayC/4Kt8oW/uofIoZezih129
H0ZSmFrZE+0d/2idp+kOaJvxSBTjMWhPVsG4esIPinB7WqFBr/nzjayRQ1ejJy4XPgNuJSBWoCHf
X5xrBMc0qvK4cowrybLG/lcm/NfTXi/VcWRjhgZPtbZXSk9KEiXn9N2C37KJBA7TWMEZrs5xEo7Y
FXp+sJBBrl1CtJ2+zCAXOAtU6k+BKGbGpCW8g07Gy0ELyH2hD5WH7+gj7o8DmkWx1FeR0sw3hHSW
1Xg0hjkHJIXTrU/PgXTtt+X8bx/lz6c2wZE64mIohqDXu+nzxVgylgtgZjHG35e4ln1q8xEbWwq5
b8TCu+LHzpO5i1qpnWebZnMzNbO4KvG3+eQuMpAuSLFIdKkicyRQcl5FH7GdsHFOhD0AnNzHziCx
8YTIAcnT5MWdSrRzl0vTweg7x10SHfjb0WrVUPKvaEVycCicj1Jne3CVkIAN7YcnkJSUqy76DCoq
4gm1WFbPHu1zmOgkrh7heY41IJcNacsc4q/s4E21HxZ3T5Xu0htZe1B1fCR14GkuY78wgOy11ujY
+5RdQBgvHRLgR7kPiS3djb4dnqx6K83NWgzQwu4hJhh7DEM0cvvVxPx8ZPCdAljCGnRgTw6cMlUt
mDXHLNg7dRcGX0udrhWLpaEgmZuyMY9lNilIragwgMVVk8IHYOZ+k0fRLAKml87PpmQMpwCU50TH
o3Vl4keYSjfQJGVONDt9oY9hQsBGZpLrrbH2xYIRu6yqeUP90x3n4lfpvxoWva9HF0AyjZSJjLIN
A0u9tHjCggpXp/BNgvN3mMI4t3fSGZhJJ3fqQ7dvPvLfheUK9vNJehpP8fk/pemX/COI5vifeEdh
jiJOBAIw8wCQhdhPeDEXz8DA/GDONpjofgUVP4OAzAV2iRGFVDqqBylnxZwBguv59M+ozRiFjTIa
zQ3yElPUH6HGJuD5+bDsPzWBPhrWep0w3MGlFdlnbQzDCJQv3U0Z5cwy/N/MQVVw5Fz7FfGcNOSp
TYYfvdwfML0OnuG7ivRHJ4H6lJ9PQQctosUKxT2LTzdTVPmKEBnCwlwLNC/LCOUis+PP93lbGaZ2
VWWadR/JEi6JG/4wYKBssOhRFjuZBKvrvBefSV7jukrEeWe38FU0gyt1NWr4nvOciCpnFe+IX8ws
zN7OU43QwTLp+vO2Yu3KkgqKM20NNF9Y4T0z9o83GXJYSATFi4G00zId4JIiVdKZW+tX0JVR6alL
L2pS2KdQo3+gpBh3UqXovQ4t6eiJ8YhnaTlXOLTlZhuqsDvpXOdH7FbApq5jXEXLnvufLNUxzDKp
hG0Znliqr079OJtHxm2N5vEsLmuYAyLHADo+50sVfusZoTw9JR9cEI2xOSHr+KS2sWoCswAIAy4T
RmIxlZ3yUwrRGFYOv6NWyptB4e+4Kt1XP5pRWu+YSGPkDrIBsz64R63mPBB9JdfixqJBzRJ8qmzr
pc+Ny/msjAJolkmIX8P+a8KblfmMA4jkbB/sVDyaBrVcXgNraiOtZfR/aLY01G+MrQxS6XRcxGLr
6lHJnxXfqBVVCFYtVTCtEznCSbi0B9ZpBlvgHsy69l+HpUOYzt9uTvmx5JuQ2vThJgayX5I3uqv2
9XXlCqTa71Rvx6bq7uNtmjBx2AOLOOKCHrGieZzG0ntxpC8velkVEHTzIBfx0R7cCU9aurRmyB5E
Sqc7Q44kjFZj5ISVUGOwfDHuKl/O+W31e/sOBOGKjWNLgN5Os9KF+BuVumYA71GYP1ykWy5Xu1TA
o5cKME9nwVWZtDfGYfKEPpV/9n1TesRKogllaQeiUbaKCs5N6IwI2CN5HPu+o+kYGhXrTHeJwKnK
EYKi0rQU69acdurA2MtmCVKaQu7ShsEudThcx5o9dBodenJ6+gDbx0BoOrJZjk0VgcUW/q0q8NHe
7dKjj0mDZgeIFtGlXLqy9Vd8vZZ92LB+RYGJG+iXVyJotx4VpkAB7AZBghkX3FBfaazvUFBiR0hV
Oqd/7hE4XDlsOZljbyTrFykgH5l5tcA1sQCXnvVSmkD/kAaUQ8gveeJIrv2r+Lf6AuZRbuFxbNpA
wbPPCuttDBdMFVVuFnPjvfZNnm6FR4Fqzq+vrEXbyNLSRfKQRorD+IagWr+MkWgQrZupP+W3S6XT
zdXs+GLj3B+PGZ4rBrX6u/tyDa8X9FTFSOFTGueH+RfwJBivdZzKcApfvFMcZ2kwi13K2JsAdBvm
Qo4DcCfAEyoohtZtMUmMBTLLJk/vkKQfHn8sQ5TOdSWU6RnfXHyF0sqjapd3QrQbmkGc+YMrV011
Co2kfb3ePX1GKISDY3wmsfazna7NhWgG9EaagqXM2X2y6qxmK3M1dxzNJvymd9hBdYrGuxxfrzz4
5nfDP5MdrSe7rte6BmsMEHWbo1rlQkziFjdm0BVqMbh08+zNRAzIPZcoeYUyPSfSGLvL0T2gkg63
n+h0nUbLJyvGnei1tg3RiuaxaIkVpXdvSlSF88JckIU2jp+pKVDqtS6ru+scP1o8xuky3YT7u6Hi
s+GlltjUxJ3cXxWkY91kGpdsEYK54Dj0OpRx75EzdHhjcMXKczeT4xpsyuIRapl7ChvlwbFJZB3X
hCfwC/It0HIbI/WVA35tB4k8S18zJgk9VoQK/c8WthV1mojyrpIBvU7GH/z+G68OnP2qE1ciJm98
Uiojuw+KRgZHmFVMUl1iSsjWBXgejAAF3rfh3ZFsGSQKACPs2KEx2TbTFKTIhqpMwDKMqdnZuPMe
k3gxntOor3o0guIggaAZt2dOtw0NRMg/5msvYorhDuX6JNmhxmgz0EOVQeCNPX6MMVhTxtExCJeQ
+RgEtp587anymgsCTwlPIgMgvSE8Jyv+MnhBCQ85CvCrYAr08eizwVvoJLWYdXnzM6fk13kajo77
zeTgTHGN1HjRBIjAnyjc9ZUTccDU+uRGNLC7/jynDGGvnqVs8zvEzrF80yxAimsV8Gu3IkQwkHEp
oIKFjOgnEATEDUbRPa5IBFoIAxm8MZ9yk8U6X2Tp2OAMeoKfGWVQHsi4P8sxU6peork3g2Y0TGZr
xR109CK5Aj0tBsgU1Z1Gt2B1OJZM40eBFh77UiIOCzanon84HwrvkYj0DTlmYk3J6qx074MltsNe
SsmGTPsAFMVhDAIskXsycl9gP9o9Zm5vPLETG3N9oe0ny0+q7i11j6KUPAHktF/brbXVcHn4EK0a
PjIe39dU+Dw3C9jxt1t3wNFCWv7bJyEaRwPmBI9uEGtJUbO7ITEpMlzs6V5R9YJa6OLFktIRyZHn
Zr9IIkq+J1tAlqqVjNPCqH10qx9pjoQ6bY8h7GrsoBUhQ9w/Rs6bbpJeesjT8W5FrqzYMv5du4Yv
qmtSxto+/ng3GJieZ+cXUieV+ysp24X/unFdt7iLpG1Ray1L7pqfVVuUUzU7czPMNHD/6ub+zz49
EZkN9W6RMze6I3384/ftwX2bYWCO/W1oOd+Sqrqym90k7FspHGnVxyyb30zjO7YggCdegUyYvzAV
sJdIZqnUCpd8+8MNkeO2OVIDp056U9C8M/wFEwmwiMdBHtufFp6aZXXxtGUTAeBl++vJsMfso6yd
S942VyQQAGcfY1TG3TeFueMB3ptvkW99hKr8fww/4A694Mj9i0tbcomQ8D7Yk/A6Cykj4mRyLr+7
R3N8rp9uASRcEbTKVLWXz6unYAWW2OiyR1LOTdyb8CUllV1MIdd+606GNZTmYRb8qT9e8LlaUnL9
4/FeAUz8dpxlyBnSqpY8XYoPY+hpJMLUces8PYjfB6Oq9uZvZ1nPFyXGv/4CKRioTkSQJLQhybP5
+11Fu9SvdhBw+BbKvLJUzDTObCWVn4CzAj4yEo57iR9OTcLCpyZDAaUzmabL1j5j1An1BECMt96t
VX7R+rjyckosPZK9npolJCMxwqeFVwxRC7hBBA44zXfZUvHsPXzDpoiHjohJUo+6B/MZg9E8rtcJ
svx6kEvC79doHy2MoTWM1ykIPyDuBKGYqpfJJ7eV0OeCDE6IlB14V5fv0hRFISb0HVJRdquHrQ1k
AMmYqpNh/+vaaVoNa8xlvAscBGdDV3f+HJALBOzn/ULYMPEyxp+tD/HZJGAh0Y1UXUWYicmvy3c8
kgWIKpwSSfm+92mO0UU4Q1Xo6zUMYCG5vALVbrIcvVmUczeJOS6nKjRNO6UPJJK4iDOQ2ziBWs+A
M1sBAjRItRtIB1K+dJco3mx9YMQFSTATQrIHW4JzImNzAmWQNxBlQNTmN/TLkv5B675iWb3Rzzhk
nV2xiRGexdTJKzYZWRggmnPARYGNk08qRZDeivuB7jugAQn2JH0YlYV9hHKRzK1cSSzseoRkdKCk
vgimJwH4kBKg0hmVfjBPG6fNs1cxhWwaX+4CwGhE/Cn7cQ3XMWwxzC7WajfdsO7GHmGMYJMmRWlK
JOGE9hdEVw7b0wYA9MILZhL6k6bZyRaNv+f0JGPZY+Q55mHPv0zQ92uaGEP8eHqMXnUT0vJbp4Ea
jw8Ip52cHb4d9NcJ/oLiuONP9OJiuCExDbN+6EC91MBBQ9K2NbLGjH2CLdOyb3ryI2DW6C9Ivikd
tQtYOXLx5f6s9qSKcDjGvnc4lnLXF8PHmODiJSpgMOHFRIDPiUJiMAQ5vGAoX7r8+ImbfZ58BEnL
Vc+cK1FYlNtUNG6CVLk0TVIuFMZPlMxZBhuKw7mhe+N/TpjCy5KybwlqVidTmJnP5Il2iEDn0u9H
mGpMs9enD/jwkABjFrsGE71XQHGBNd/SOMNluLfnuJRXyZuxRJIx24nzVys2druzNnRitXb/wL/V
MVxYWztmgswGul3jzXD4mzFLfF5NpKEov8zal1N8aqf40tq8BTbrpJiIAzw+jx1hlZ+FN+YT9Y2T
VxoLi9jzuRkXhMNBIicr6BiwudsKVnMHbgEy3OUySIKloJfSeBpmejXW59fB6B07lkgzMGrqfCCk
bbZHZFsyWeJ7+Vv0B+0wbA7GDS6hi9pQMligd91dTt4Xh6Nd/WjHQpO2MCdV5KMk4pns/YFdimBN
D/6agks9gPifKUwRB0nslqlnQoVwFhgf/itU+K976X7uT2Kbb5WzoouMt0u10R7XyaDzpzRyAYzD
tZ2gn5Xb7EGMpDXUelg1M4iaEHjK3pvsRWmBCPsPRNrVMZiGIVsr/VNK4E++tbAhZ+/UjpzBc5Ok
UiTVrQD5R8GGic9n6aes2aWwRup1iNVyVOYvnXaW/gZm4l9QkGkWmtupeIxDzE1GjjjC93WZbqB3
iEFozFYh6PMPOY8C85dmOgWEdSOtBUjgeE1wdwNP7M6BZ8TQZFZGYMNCG4f68itYOirqwLO9/k7D
Dgk4sd5r73xmxEzMuPxlJN2PdoPFsfyylNs7H7gPCBD/RKNZHxjZ+mbzIaPWe86CwCCFf1mmHdZ/
uRE9nBy2GOgRtKKpqsAs7WydarLUv6ZTgYVbCwig5+FhhFAn1pqUrBPSfr6UhShFH0iVJiKGvrfr
CpqdSabNYrgHlx/A7S+ZQIU+CIZOfy+gFV4KqzHtxzZT4YtZOw2b7cZemOf6Fc9Ij08ZKUgW5CcE
rrBlwK0qn0wlGmMugf5O9KPMhVGEhy3MKGXKo4AWAHUJK9Ye2WvGDl93KRqXS7UoYlPQVsmWf7Wj
rjN+rSChQCLnL6lsmkv/4MQjQ/8J6QdD64V4f6y78bM1vJAVTzmyK6ygLcsPifkOXsHRXgA24v+L
E1k9JvzTzfmPgxGIUTnJoeJqU/uiFZijUUkRcXfT/GjwCCjnjwIXgHm1rmSw6P+ghaAzt2uDTeGE
kLflv6aIOQd2mIBl5jbQIIl8WsaRs+/NgOWBj7z6zs3pbH6At2UaQo1vxiit8SUrusiJbojERsp1
WkDN0IkXOwasFtOxm5HTPyPgMpIooyIyqS2cooIKmwSPAbh+vvdBCTn/AUODYXJkln0839l7W0Gx
ru1wMKrkZYEneERs6G8NRukbr5ykFVlCPbtOScB4DtYJgNbI9pGmm1wTCcLdMwbr5mYzSLviJ6ZI
ftjpQQ3VpAONDW49E6adXAl9FCPrdNnTYslhilCh7pY7rY4wlD2BKOI3asadO/csRauY4qMpHeiw
oNVezsbg8Taz5JhaeKfjh932f/vlwc6CfpOSlxn3L9K6wTQK4wswfSFypFCUfhAtx318aAUwKQOL
HEsjlBMdgOWBsCAWCr5zM9ZSAfFFsecGVSHzNkyr5YN+vISblRcVkDIbmCr231GEJRhKIys8j+Fg
RVBGor3JhZ/w3xn1Jc789/LiNbU7fyDmGiIrCFJ99Ea2C4lXUaJIXoKazys8TRmaWnI5g9BeEcja
fmk4aaf1Api1fDgrU2KS7Fu7CARD+Km9Bli5bOSbYnFzBPt9iuR6V+I+ksagYlp5HonPciiRj3hs
EcpQsnRaICzK1TPE/w3PBbx33ahpXnkDH8plXWxNjTZMTphUWoripIuXm/00d4t3We6X65nDccls
7ubKme7/b973T0fs0Dbv6C4dxTDut7rZSU4zQejPy7T7chKWbmf9RQc+6YgobVd2nQs1LGI9LENU
iXN2CGO+QNczyXuR6qbWGFUfMVq7/zDNVP59Q6SQwhZ/fsGQglpYB5CtdaqY6zohZSwVz2dYLC2E
zGCK3SC9ZPP1vAdCoM3KPyBLmEQue0bU6l9xdNOihFD+08l8MyJBRai6UMGd0T91dEOzy4tv36eQ
9/8GxV2IDtyEV1AJ+CnYGXVPIkDgjyYo195HC2w/OstgzVQVenMhIhLma3bBMD7fn70zYozIMbML
tWxQCte2WauLGJUM56t0mgVhDXQFc10zA8Huuv7N4o/YkEbunmGN0psPFKJxU9YYzN429KyuC21n
k3fzw8UXa//PvR7TID1UWQNcjwUr77V3xEQcatPcZpwXDqvYGEWnq0gO/0rr6zsapeki1wcKU/Ix
+OKRuKsQdboqH6R/rgJfDtU90Bv0QUUXQbKVUOFtXWXrLQB0vHtaTb8t/5JknETzz2RoroqSUjXy
65Lfjrv2Tz70p30cDH6vEK0evi8pyXCQeLHjht1uZdqeW+6uvObUjTigsNmMdljTM2iQj9wDjFHW
FxQDcch3AUBTCODU9dS9W8giMJ+iEgGhfj7oG+Ep8RPBwUWJSjKEZ0lEi3wA8NU26NA64eQquC6h
KU883Tr0Lem+uIs0AYK1SYi1j/w6i87qVFQ77SVPBwYcd0LYBzNL0OKwjsXO7lM+MgzVxiQC5wzi
eT62jeUZ/W3BGooX0q0uV8+XECCnJzrgXhUwFscEdyC3HN6hIst0JBqFIH9E0fySTZKo/6vrOaJP
+lKoQGSWzt7etvu9tM6BW5OPPcVUSZ/ffEgOqwVYlGbBdzkfa+aOpFAYVo7FjiHZf2RS5kIGJaKw
70Jz1wsG9HBgv2jCmC61bCNSBWZeGxPmyNKd9CiCZYLtq2/WiekZzjy49vTQzbIkjE+Wfl+oHasB
w/imtjBdViYrWosrb81Qwffu/IwQ6MqShc6DGmjcL95SZB2tcQ/xB8ry0N+juukEQiF+/Ktmwvhn
uRG4bPAbWyMa7ae5dqK5bfGaIOH9iD6KYO2HR2A18WlRBE7Rigxmu+KgxVULqTMsWVnaj852+oe3
VShB1xaSGmiKvkmFHmu0i/dkn2BelRsHH8sjEHbxBRkJRXrjcm21aehIHL5ZAnDydnRyYub95tFa
8yvpO2kCmbf/M0+ZMM8nCB9cbZa+7mFbXLI6VQ38z+33GVn/+iwHod/9ADVE6m06y16RSt+St7YR
G/YEcKwWkgBsEFOhHG/yNJ0xOjPfYoa7i5RChePn2a7WK1DZ8RgI/SqBjazMB0KoTNsgEAUlk3zd
fWSy37vjhm8HTW1N8YR0q3EB7YlHrjiE8ol5EnlqzziavCPi87T+RoDzOypdmGurezYWxG08c0mN
4zQ2K71J0MqsoJCXnb6aqO8mIxIfvhtbYO7Cz2ASOEnASjX0ckrNVphugaQZ3YaqMz/MXT2wP47b
uq74aT7uR+9mQtHcvn3PeTAHJY8qAkjoMU0ztKEe8pLw21Bnw/6ThU2eQ9TEHKYOg9U0O/PfRuf2
t24xJmF4seM3Vig5GDm836Q59tNGSPZxTMWafvQGCSIaCIe672ozZabWNAuXXxMRWOpbMhMGi6Ps
wQnUgbPQn5YNqaMQBbmV1a50vAzpOD+Z0XUrpc//wTJJUj1ceRKGKYVEJwCuL2vV1BiHE2yLmyKX
9fjA5+xVbQPP1xObq60rMg3QUt98XisU80/Pd+2dyX/XbWG4Y33L021bhVXEcHPQpJKHCnVGAgVO
a+izuhWADBvQS+wpTab+NovggZsPKQ2LiTlOQgHD98AUUH/ko41POeXgLC3LYXpbrlk7CcQ18Yjy
3UP7VsWHRNSYV3pQsocoEs4e+8Y4ZsxWfT6kKSdXCtEAIETYryT52G63QUnX88ddvTknXBGJ0/t/
DERfRjEKHaIm49tpTfBlX+teC7vMWYSRaJ/loKjUJ30I+cTopulW5eN6FrCxwE4NilJ0k/tI57DV
F+DIo3cgfrDhW3nl8GtbHNDr8JVIpWIYLviQkefJYlp8b3vttax0yebwBCyOHe2/vaYOUWFLgaFR
jEqq9LenzYvmgfMpb0Hlzf7oLe0ozifo8bgU7HjcAeU81/jQgPXP7ZmfczszpVKwbEv2efTmR616
jfbSYmnkweZ2hSD1DfaV+YdG6bUwRjk2dEasjYrVFhe/1urvmjk1PGoYnRLaAbEVSx3y9oP2ATQq
8pkMTSiIplzAATeoGIEAsypZQeosSRj+5mfXolPaQni2wSoGPpSpaheNPAaXviGQoYJK91n/CspN
NgWx83ugOCE46DMkD8lFeVLO6WLdLKwVC2v0EQUg8oKyvZ8J1zYqfQ8o25/7ftSOmj64J0DpDiEk
uTPIkX404dH5nqT6lwdT+9Hz5P3mzwqnfFU9/0y0GLDnMndKg16D1AtsdIboCGH9tYWYMpkduh8N
eC6VREd3iGI3/5GHv5z3HL+JSf7gmssPwzhBXCUH9BesKlm5+ehRmFOJsui8DsWwy6YBkpANLJZF
wo+LQWZJN5iYz0nf2Y512+W9F+wI0fcWrObfdjPcWjTFQ96x1SJFtG7tAmTDZ7DVhJS/eeHItO/s
m3xz7OVdYjWJBEiVL8kIYXLOtlvpES5Ec4Q7hnMD+cPC4k6/aWX9dkp+YQD+3bYnygo+d7hbQ0iF
vlZ0gmnZox+Fo1x34V20uijS+ANjDJilfl8vvhk/izbFWQJG7GkGvisMVrUpsEiWQwU3UT+3ORLT
29jQIW8lnSY5BW344zHGB2Fvn4fLT+U0wDy/73dEZWCb7pmG9q0sYSjUV0DZ/jMi1fIElIBa4k97
YLAxKu2aWJihLtgh72CtHfSBl8kdxqSaF5433qtFLG+U2A2TQxMzKwuVWTu6IQS3h97aFavWhU9i
g+HpzbcULGY6d/cFBBlFAgwbiRf+erXoyhRVvVtFtoUaHMplavRzYxYSwdEKi6k+cvx2LLHg0701
QPGBwqmW7YTOkD9HOdMvwdM0wcNDvTGecDy6FuBC9K63LFYJZ478gu6/Hgyugy7Lpd64oOq8H3cz
foZOs6B2istR/qRfXYXF0eH/Vg6T6zpHzBx+IxrlQU6Lfe2ySJTNnpZyN5gIdG3znk7aLY9E/hEh
DbpdyMGgkjVBW4OxPDRRBtXt9Wx0r52quPX9V+xwblquHxb9UcgPusWh685s6UK63vxJJsVlVlYw
xlVXYAPn6lvWQRKonh6SH0pBCRW+DKidDUdxwB/yqI1geYo5RKWMfq3BmVjqxPIaL/Oe/ZF+2V7V
xHys7mu6k+UR80RomAef++umiNsgjmD1WHzOyPfmeuaHPxlHCX8AX4GOajg+6ZmWKkDKBjM4ML9W
OjYGxA4+kAndE1A1CpwZPVtqlxqAzl0mzpU1GCTdrssP0dIctXsF8UQ2233r4FSRSRGmZH7YHkAE
SLajsW63HQOnGydRzPoIy5Pr6DXaa8I7bM2vaAqe/tI0cjUjMLyU9rPHa07DKCSwHZ87hpuHi9so
9OsJqusjUkv6lCXjI+a7i52g+rqcHGrHg7ObZ4C57b9qBsNpcRe36o33eWSU1aEfxNFVlBZlcky/
tBL4IeKi2P7xkULDZfFtYz4TEiTgs+Lhu+UgiMTOYhs4qOEgAy489OwyUe4vHplsnPyiCEm0KTwV
gf1J741I/sxlbNZdDRhHS+xPx7HcgOCEnDqhP+vMVs4ZC1uPQVbxJwlTU6X/gLdM18mv5fP0s4hO
gg7vojDAHfM+W5TaroYlUw+3ynzOsjpdWzrzS9r0RrJxQmUMPZwZgb5Ae3h8sn2cwH+yaHGIbfza
4ckvB/i4jEtd6WMItTPEknQ2OdOyHr3o2QD0VEFVLz51uQuvToBH5Gczb8vRt+pj5uoGDGKa3P6q
ILABdLovt+UGyb8XpJnePARcBDrwePYQzgYd9Jo459pYElv+MbNWNjQQRinLtFrsvWs+CoPqB7SK
L8LhQ/lz63FeDtrb+3gvXuVv9D35N0RX644ybL7AN6GV3IjGkOzaNm1xw6QGZ39ML9yvNKTJUTxO
vXeiIJ5LhnRzwT6EVg+vmhUw0QG6PIMNc6uAWierTsUKDQrrNGfQCWy+ckECDePSx5I4FpJAMmdl
mzEMjrbwwnzmpAe2J47vDr+manKN+9vBA+XruSkQIH1JqRCuKuk44D9OB53914iGoks63wnsdZUg
uPa1z9M9Ft0Oe+pWWByrVoAjkIK7Osgb78Ge1/0NYmLSs5PsfmOL1+7+utqdGxVgLeA3ukF/mOa7
FoH3ysCWIz0CMD0AhLOvbYFtUldooyV3YjetOLLRevWZgXAyxUr+IWvvVC68yQoZumvlBOEu5B+f
PGf9oa2n1FHjsajKSQqqgBXaKk3WIUJD6S2WQ/LKigIzgkRVbYKgPcPkR7+fHLtwNG/KoSM98zMU
NEEMU5pgyRkEJRkkLRNycM6+Qb7M3wDpbKLuMTghgj0yKHecS1zjh4TuJJdQUx/luykQSYEJiuYa
bYApaFoyaIblu3gsYno/Z+mLZ+a324ASbRiOD3BGOCn9sbvw/q5YI/V7Kw6QsreXg+EOVetdCXRz
d4xj25sIcnW3P4+04ylb/fpgMUMHeBI9gDPCjen30Papl81C9h3hwvfnnm6UQQLC7MP+LGVGRKTq
TRT6oZW7EmfsvzoiL08ct6ssSIOtGUNdCNUx2fmYu4HD+ScQ0/UgRfA5tih+bgPULr9P5fJq8sbK
qZpOUu0m8HXxRHk8W//ZT7topaBWAMFW64sltOdWyUh3kuJnhYxoWayoxpl6NCab25Ecn53EnIhq
nczaSQ6Qqpnzsz4YhNNCwNEpcQCkUcAWW8WIKoBtREhVhjkMduurGukGSR+dE09AjS5bLtAyllQR
bv7rVclcUBV8mAO1jHWhzU7BcgAYkdTSvkJQ/3jONu/Xr5fgvsKDszBG5EtymX7xzpGfoYS/6Fqr
WjZ22fsPeE48aOMuNPmFO9v1Yh7CahcDiwGsyHphER79JlJKlUxXBkYmL1gaFRTp4J26ZAYcxWWK
eLcUdU25Stmg/I0dQvb4jPAV8Sm5AveVLKNMnZFef7s+cH8i7YYhhRhqPTsIhw60UAYJmuGmGhz9
lTfUGMNtr/BdeQTquP0NE3FkpDx4cwuan2Z9NT2sNDt2PIWigWVNOOWJXWVdpR3Qs1c8RnsLpGYa
bxCqWT+osHz6b66MZSqsmz+ek5l786wWTZK/jXGKZGmE2EQc67vXx+fGD0504h1M2X9i3uyx6FXo
HYGVxweUJD+fePkZmBUpAgzvw719pEGisE+kdoxQZBMMViixOyhiCPvr9B6YZALE+06iJ/9E3QRJ
EfJg7idQ0P/PXjZS7EvK4HJxbhVDq7kIt3g1EkcyMTVYHJFL1cYbB7NaYryuM18w6xRqltnIL1AI
gQKXd/qLsNa6P8vxH0JKs5U9TUkL1XerXe/dusSBP5Y7iLRshaKvH58b96CaB7oTDesm1o2ELOfY
fMUJ0n2LNP0t+T2aiDMO5fWosfY2AQmFRFC5e8nEBxDGdu2f5AMh8MdIiKTJRFNf2jdQLnuxlUdx
Td2zZTx3f6XYXPi9z9831ZmmC91sWNexWfdYnGrRV4sy1/rbqxDxPYg/+4vS+mq39CgjDBMHRl9O
A2a9R0Hc0lvW67EnRjVxYdnk6N77QG7vOgsVQGQ4X8S1mK0AF/Q+0FZzomFcqCkGoGfu8Wo6/WgQ
4cOpjmt5dO9DcXWL3diIYe3SzZwQY+zlTT8vu/d5m/3rz/M6JXBUYIkfKyPyVQbC+E/eMLgXWaTH
uXHPxasrqNKwoEMz34xq53tH8+zuWOXwhsXPAL/bIi0sLq9PABu0hEE9ijJJxGtB8XLWkQuTJxx7
E5yrqXGzsQdvadIh38I8XKeXkwVg8Chx2dIpZzOsdh537QqtgCjfIIbRsmRSwIPzEecKtySHwGbm
CPoeeO8ybHWAkSgcS+CyjVZ6yPkQrzVoQKLU/40+5B5is50N0UFIb8Su4Fqb9hNcH6OIbNoBw76C
YZkMFf5lc3T/oYiC9T0wbinJTLElZUv08eHHPJno8nSVTJvHBkZ+R6KfmMIpsAXfuThbHK8ESVWa
mgunPT5oBFZ9jAtOGjCYh8Qq1/q4hFnm7BhCa2uq6XUvoWMUTkN7hAYEPVjwD6lVcUgJD8xLeSGx
IjNETyqw/sTfYykDqSsJtl3QaiTxBuX8nX9lm5RJrNPEMWyezdjTHSnTEmoK3KujEkdr9avUZ54V
L8N5jjYd+bAZgNUzve5bsu45YcTD7AxHgJVxehyqQ4tQkpXb/S6rY8+15iLN9UJt4sNnfIKUwesv
LgD5BdHpgmjN7vT3PFjz8+q10klM+qhL7CkTCmJT0uX2SERe5swmVhsPqTd2d3G/fdSvRxpZ9XXl
6MIHmheUGnlkSX7IWEphC1FPJfVgIdRzcBClJfNXhWUgpzPAl3Mp80DdS1zlFU7P0k2BaKG9k85E
V2K+ZqUb+aarWlpWxzlvfqPUQyjJifIyCS8clw15fNuPiKcaIsD1WtZize1VEbphnkUGIElrP4+e
iFWj27vnpqWEcUaT/PR1XT+m2l2wHsFhCj5ZT4n7SCOty9WlCl13ibvzfRueR5b1FwrrWitomaJK
8/1bG8Jb+zemyGhTJNQV5+P9zITd7rm2+a3InqdZ8tkfyVP57tI4vbk9gUkNYOK0g71b2FO0idOP
Vn8V8PedZV7GMM0+ICgHzAdCQxZ9n/BYqgxgOrd/7H4f0bSHd1ON/7Owb+tYFxMaXUgFVQtT7V7E
NF12cyfVBmw0o8wxoVVU8BcIn70bhskhrnZIdyBqjgpPEGcrc8UfOmmA/YYM3QQ5HGIi+ggtI67E
ecZEysdMCAAiVA4R+dL3IFVhRcSqZgLBpM9zqHJkZlXnyTS66B6DGlkbRmG+l0EBb0A0FnhiowbJ
Z5mXDMvWeMYBy8OlwqVO0tS04eH+JZQQF/pMMbH/x+N8rK57n9+p+fL5LHFo/tOQ5294IN8ZE8HK
15xo26SVM662PBO0GUIByzAEYXe2w+Yv4Xt8S9p+I7+ZMgfQsKn3wd8Lfxo5E1K+RPE1T0tlg++9
joHZQHePjlbkHu+nV6dnHl48SKSfiqHj8+xNHc0evOv0Z5o9pJAdFSWROdhUHKmEwBMiUTC5FqLv
TYtnLcD72Iba5OC8C7lNjR4ANuPKS5UoF5D+xLuxW5VGGIWaumGzWJeNSccIAVhRmCSfrOmaiBna
WjeFuXIMImkxvcpdWW9VT/+Br+DxbawZ0p6vzyfWpPmPW4LYrMlDKS8uR9ZFIXhPKTFjGgPKiI8L
oXpLpvtVL6BxOj6aOw2oKUFZ4reQ2TyxredsnZAFFkDtj8PoZhyV2LmZRm7zpW+WnwgCQRaNa+eM
MmAy8fncbhGkNGzBudU/Tl/6S+V82q6lnnTXXwqqhxgT6UxY68gNY5BvXAViTYwltz99QYudaJQh
fS+ZZ1riT7O99dPJm9V56a2rmHUfh7Du4x4VFKrtWAbjmm5wnWbIpl1vz0Rt0OEzUgbUUXmpdJr5
qU7UCAdGdeH2rSocX0WP5msv+gW5FAmRRX7tcmu6ZiHQEzKrN8C1ZsMKN1y2yuTZ4kB6g6YzjA4D
fMQY2kt/+WkfAKqXMGNUOxqeqr0dAzsY/UoZzYpU9iuZ067mPWgOTFqIp9kvQjBIPxd6uZzesYFI
9egnMQPKg0Jq7QkoSbyPDEmF/Y/oeLZc6KPHTFnI/6LdOaUSHS9xL0V7RYT3meG40K9VbsQFN1ul
G0u3ME0QpeGWdY9ZVsoCwuQeYkoR6j5Bxi7I+0fP09440LHq1mAv2RymH8X2k3NV6bE81IL4q0l6
c1mmJYNHLQoOft11BTzTHqvlPfO6CCH1SUsuPXnX7DuRZgACfAhfFgL/CYzg85AxIFSRtS/XuD5O
aglivLWjSEJKlg8zEdFwmspfYVA3FFxRZJUDcu2PRBeZyxqjIiDTMSBUFVRfLVbOwPuTKj12/tVx
/LKNlJzBQV/6XthWmMNbuhvttDfnnqvQLW38Ig7J94NAaIox1/z05/AgXfKufZnx4eKr5qFO0rzu
TA/q7UeCs1QOb+ChXwFLfEehQnh2V4G1z1tcukkzcd1nml/sSSalwbj8Ngi/saz9KlhQNPzN3Z6c
iWwIlKQHPKB3gPdc6f66xJWXkzdeDyge48yaaQzlEDx1FxGstIF+5gvTH5CsPQyeuN59Xbcd/WCv
fx2jSMaxCb+L+Ro7K0nN0jUOF70KgFDf9WIqDk2iz9RQ/WmNZYFIyLe5WeS3kxc9kOuYyKoCDukO
P+jOcF2hFAI2yyJCB7mww8LuOf/zCZQ9WyI9OKQxuY5wqbBT3CkT/WLIIzHrF4FOvVxJIyLqNYbD
VQPqv2oEUcJoxIP1UM3J4NlXnGO2huw9jv7DFyXDCX+jQ5DqpIk0Y4ELmE7DkJWmyN28Im3K1lGR
BetzFk+AryTp7XSkz+4YM5qc8NWB3C8/RWYuXik571LA6LmMh/DpMidJxGdqMSVEe/xc7Jag8CM6
gtAwyB+oNWKAHprdiWYNuiNsdGsvlp6qCUOXXY2HaFFotEoSmFQ1TP4kKZ70qFsCWzUEZqU9XmjS
kJ1MPhJy2kQogEKi3bbLcIzMVlYLRMqyCOF1NAyURKyjModQ5nOVxKeBYnyie/F0SnaD3OhYTvOb
ICFK8hgazvq7nHVYCc0teAhPI1xZBYnG9adBvQhy+qTe822HgqNczbAwmcqOK63sZN7MYclTa07+
0o1SrIoh6dNStHINiyXLZIJ7RXG/ka/a90D9nAD3l3mimjsFbfPOuFCkRn5qskuC0bROKMh8ZUcb
vrkNrHpp7GDJkUGI0vEV3OgJNHtuwBfMkOwE4gYF9j/RTnppOsfO5nPnxmbJnk9tBP1XsJ+YX3VV
akOo/iZ3a3qPeRzLHWAS4D4jLyMKseYKYgNxzFI7kh+sU4xFdhb0oi4Eeb/AWxCCtUDbxpGOm5Z1
fNvrPx6/qtGVKeU5Sz84HgmAfTGUtxahWWUhy9nH1q+cIDmToZjXfo3a8wUGp0uCmcEqcy8ffC6s
UP6cQPewxpBM0bG3/mXcgcijcSNHFsKQF5yQb5XnAkaBYyPaSXZrXoE95JxX9fYYlDEAKUsGgK8E
NNReYxF+B9qe3b5QK5W5zZl/5him6V7sGss09StBZHBotA0NcJvva6hCAtFV6Ll1Ro4JO7dyHaS0
afbWkQb+vEkUP7zsmjOj/ZKlNWm4fGAg8p9UNH7916zOqxjJD0mVR6BMDgtn2EuyWOs75d7ZLR1W
YkXA8KaAZYUW0v0Vfu5at6kz6E/3lq5vUMZ7PN0GPSaytpG32mbW3mzt+ilVMZIZoE0nJUmJqk7I
54jg1kwHxugFzPgpO/aC6kN1Ih6sjUitYbGBfaAv9v8SrrHMc8qaLmfe6ExfeJIfJJOQazTpA8gX
kGxHp/1K9U/n62sy5Y9B4KjFVaVs9WjOv2ORVCuTRDLp0MSJ7XHYn5fAO9/awEhgdvdnrQjR30AJ
eYk7FL6RiiJFzIPWQK/U6xtOj9uOANn7lBwcV8BV/pHbNRx+h4cLMaeAar4+fSrlAra/rPdpwoJg
KnERjmcNhF3ZJAvvcL2t3gzyJ1LHNzUNS9jrzUODQCNZp6YZU7zQrPPTVmXe5IJ3ChH/cdwKDEvK
dlNBpFG/rrAyJI4Nh9ac7tVBZsnZV3yqMVv1rfzNWzRBqhNIXX2qYqRJ2aKthD3CXLTeTL8hGlTF
OXNHojhSIBiM5ASphajZ1MymSnRRWbLsbBF6JMPZiKLHpVvYvnMTeogvdd/o+gO2kNjCpEloAukY
3Z4PxcCTZJkvG2n7bdKTvspkmU2ZgJQTsJu//adjNf1eO60YXD4ULL0Og5bs9dEu4spBt5IjAD8w
4XgTv7I5y3OxwNs7xRQz24T/hQJegb12qMPqQRsIFUlmMpQ6EQUPwtFtmLo/5jxFKDjPz+tqX8U0
M3ljpWoWltJXeyvQLl0Z2Hvt7spP9Dr4v3pdiLIMrLu7cz0lFj75fpkjVUZeXd3r7R2rTngJnjru
t9fvuKFZb0YYTrF/Ipptme6boqNBj9s0TexKHW3KbQKeeR9Ly4UiCwO/6hq6hOilyp6b5ivQv7/7
guw2jfXmfCrn+5SHdgLeYsvzE6prge5qWHTb4UaQ3eq5Nch6rRKswpMCDvkZlzpZ9Qxm4JY8MEQL
Ur3eP0Q1dQlFCdmG1rbJrO8ctw+nRAq12615DOOMcPrOqnax3s4+cbM3DcpQRz6a0L3U0pKeuMf8
tXJ7vh8efyTOlFeF/q0b/k9/Py4OaZZRtUvxYZkdE1Hz+KGO9O525VFJir4+KkV5ONuTIhpKi9oB
hoy7x2Goht1Dm5m0WxDAUtKF6ddJsqjt/sl4orYQ/I2d56VTVAgdLX/Eu0jCztOry338xZa3jUEx
ncWBKzKXIe3MUmoGgWvLZcpFkaGn8pW/o6rKlH0i3LiWkc1LKcqTseoS7/QS4zC9GNWeuXIHqwQ4
OiLDk7dsqF2cxoRPswo26VgNwvxn0KTAVg2aT73U7oUMq1aehq/FxwuSRBU+m/jXNEsz9vuB6slX
jbOp4iciUL50Etjd3+JczPAsksCBtiK2Y7icstg7ozFU9SRj2wa6F7jJhfjunUsJ2pFIX/eOtgGE
hV8DeuWKmSN2PoA2erDw0IKIuwYjvAkX8aB9VnSJNaiSxn+wUJgS/q4uTr0+OhBP/2L0CC0s6AmB
rI0o7QXV9M6ENwiE4qFCMXdYA3WuCmNiFuZLiDdTa08HknGEe9vgzI9dSK6HiEOWCNlLXWC1Qwvy
bDBrJpKXHO66QiFYIw74gRvnJ/qvyLjNLbkWVToAvmcRCnFi/OsJ43s9Dw4rleZs0b90d0RNb6do
rPcBFKDVRAoN3mc0OpCvngPM8rExKOmqgqEsbTlmAaTAtQg9vlJnXc+W0DgjOxaK/T49RjM6Rk/g
jc65SQnvNNFwCw44h/8rmzf3uji/mZ6CxNvC2w7QnRKNXAWwcpS4LQdbgybLi7A6iGhP+S4XM+F7
KWOjJ49+Ai/SlO6KgaqTloTvfRLsEzvk241Pt1yGpt63vyronpS88ZigNQkXFuSAIIVlWDbM9DW7
yfePsjpnsp8voJy+tXL6G6XOyBExYoeD2Y5Q5HCuvAvnxG9ln8l5wZzue0NGJMVnWu88CfhMCjl5
XMI13JLs+mPn7TGx6ncK0XFscFOQWwP6wlnfixxaavtn8O+tm9Fuz4Ewb/OoapeIbhnoiOmPdIGG
j3QBFhku6l4bCNJ5Cprp0ZZNTI8mqhW1ePdVCsEzN/1uKqq9EoiPWb7GOwXvYJPnhX+Kw1rPogYb
vqF3SWIRf75xJkaguydoghrCWUMZ0bx0ziJCZPoK7eOeo/VUahOnnXGdXUNaaNYS4xqEhk99L3U4
NqOZWOh1fO4DPuaji4VQ6u8eV5TLz1w/7a1mC3XYhF/ISqgJGGOfS8ejQZinkW2LWySEB0QsePwA
7oUO0b1YVJdrXGBjBVna9SCGJrtvKzsaeNaM81+AC3CuxKyEgh9M2UuVRSPflQJAS/D/UjcM++lw
/NB67Ieyt8/OgZDAGQqw/2vSNERpUsASR2LqyASZyTIqHHkPmPaRA2MDPpa4TzqesBrIQL635jyv
ltyLX/ECNeJQ6cHbrrjC8ENeOGqUZYKCg8qlIZuyrRIAkwQimDnJl7ScZ8hSs0FcymrLuP3RpscG
bnZDqC8OMzEc0guaNLL9XaxcJdvSkqKAWy28AzaEDDUzfY1nRNt+/qm7qcbXHjRwCyARBBdpfTn4
XdoCByO8Et5Da0RFi20U/hIv/Cu2UNLjomDhlkiQ+URLkgZIVSREcEa/gbeplr6Wn5YpPxGQik+k
7UJwzRg63bCsCvtUtR4h9kUKBKr5TNqMQe4T/9iZuY8cj8EpQbQBTrqp/Jexwhtb8eAJkTMlWO2l
SXLI75/Hp4Bh7iHTIHHr7XaAGwRgk8ORk9tslyQanoF37z57BTaSP7OyTWMFWOvPFiaw9inXX4bz
ZdvSp50WFjenlvueGlrPD6giSpBEIf+a0ALBVMUAXpPjfDTop61rxNRIjE7MTJmxW5ovLN1doAvy
mlexCIbI9rMlWVV4gpflNQfGCpnoU/Bi/DvUT/NDoF7ofQOecFDopagibKCsV5Xi8OdHh8j9t6mr
AAe12aIT6vGv2ZMFyrXPCq9imZleUsEsUdbt+nR597vdTe/5wa9fvwjGSgILIBMDvXCVqRNHoTxg
nqsl3LfskVk4BaiUG8HgEuvP4NgJm79jKOvTSS9MqTaBCF3B7aegNGG7aEeX0NmOlSoohQMmkT37
42ggsanfTfz0ATOGlmfp03LoTd+U09TfGCJUPRLCKOogZap8VV4z55Wk53RX1zC0z0lYfjBQQn5y
s09V/p42rDfBH9wViRZC++5DVWe8QgeO4lVp+CByoHj7/Zi7ZnOY7ayKynDL1r19dyHA9wio07Uo
CRKJsKDrTtD8aYIB7VNBKnKw/pVVEAIeKrwuKREd5wB7keiMtIM8BTb5SeRGmo52FKcLnCctWK/q
j5tPz9nBUQYV8jC0Fu2AbyuVhlc7kKMRyHItdNvEKseB4I9Upqcif9/vu9qTYLdOxbzbIjhOCuWP
aN1BkQseE2RDDx1Hs1al73iRL2LGSm4q8nJ//c5MiktHPLqXVZHj3VxlS6+4Z8fUiP+WTgqxwH8E
UqUgcwsBGRMN1aCguDC7wYQiE95+UoV7zf1QatFRQaTv14/kx3P9337Q1xJBrbRoWDz+XnfdPT2C
D3w+MqpXMau6cVv+64VFjlRnDieQc47IxNAO1LalxiInmrAZgDkEZGRXVeEw7PZW3E8JVIobFaTH
y3rm/Dsbb+6wQv7F53Q8xpWsepD8uNsL20Pp3q0hPSjigEhYHoA9A/BmLWo3vYv7974oSG2GiNYO
dS4F+iE3YV6hF5RLla7/Gn2NIl2t1aAuaS6goSxMP8GNjEbQEXuWUuO6H1tk4dppiLNht/J7S7EM
S7eaSf4BGALsKnhv5+4s93zZPse4NBsrCPrimh8AJZOysWmfT4U9n2GVkAEaYkxiyQhpcHb0gexl
UBnktzSuafCwzEAKGsPYRM13c7VXhhDCrbSKzfKXpVYgL5+nnGGZBqTzdweG6ZPU6YyoJ89C7DyO
HljYMnpoMaxtJPzLAkcwx4it9yUvE0v1gD+V2X47ANCehZjaEz1ghJxuFXBxQQqp83isuwRzeuCB
uAYawKgR3oupXdfY0zASRVrJY5BwxUyXht6pOwIvVbErGbSHJQUthO+4k0FV9CSbkcwiZwjpeVh2
i2wtjm5U2elqlV7dLVqK44rQLTPphaGEdtb6YNRw5Yudh10xGKL3vm8dHmTO1uz3BakWaPh9H7BD
d0QzKjjp+ASG7GMjTZDGe/saVCLc5oFMoLCZaXg5MxHkVUQWxDu60KcEsvEqRAOFdAHEVGFVQ763
Ha4HpVl6icyYf0aoKWBLPrw9uWmvjWJPlQ5GzzflMM45BfwhvyQq2lYqJGO0WFjkbCX1xZF/uT0b
Iy68ADXDcatBr4KtN1ONj/976zUTrFRwrkucPBvUL/i/YbsbxRXARp1AfX5iWdVNmD+EWYpZpxZ/
O1qQee7L34OdD7H5L30Zuk/ovBg8JfCfoREgy1u8z6pz8ATfDjThlfdmwAsn8HHRB+G/A3qOppRu
Pjxm0fzNbHHZ3GhHFeW8Q4Fy2uj8HeFei32dQtX/df93J6l1DcxAfhnsQ4gRP3Go6/4xoO0I0f88
1iZltZiRCNlg8u0DTaszcWOXeQC6IesnD7m44u4EqZMRWfjmHNJDFTU8qkEPmKBGMBZS1+XPKKFm
D5ypcDS84ErZxXyru6z5/mqqNkEGQHy8a0Y0ueuF2GUdfIMVy7N1bafONUhBlz23KpXv/qDp7aAm
ZWndK93LDknpXff0rG8xWtZy6TO1/vgXTxGe3H19h1h3sTuP3fEpJr4H8zzilBruYNaEjFW4Sh2J
rEXpJ+kOovnLbGNaBOWfUT188RCMUG5I6h3BNnrqNTc/YTP2u43O5a9lO0kz2pwMMT1L5UyGbxTK
tep4klCYh0tDDI+IPWD+aJ0SiPopqHhS8HlGDbbsDBmzDhurTOcMhwgDlH/j78ZhhKGKMIXqMBLt
Vh09lVqOk0zLDedPRdV0xhPuVXTaoTlFTMY79hcp/kbU7lTDjAYwSMLd3Flc7pCVsAol9c5M1xbF
njVqiNyohIRe0Fs7YTnXtqKUtmb6Rjttx6sK3vphoc9lO4FuUY/X/AYSaqNEpL0qcCJPbW3zQIFh
HKdPFSMZ7jxMT5Ze5VKGOAdtN7sUDPq1Yw9WKo6vfEL2Q9MbzmEYF15UpCUZ45QUoYFpMFQavneF
yTUXiv+Fbm95xegRSeiFRZo+fe0mTH1Qs4Jh665L8JMg4BF0sBx5wD58dsYtZFygI7zdfE5dXVnf
u9KW5Ig4kE506/I96nIAg9IQY7SOrifE9t91HpJ1Yfz263c49tAFzgTa0nixuJwSk/JEnpM3678i
sHAjty/TMJve4IUjq6HXJDH8uNxE4zFwlU79fYyEi1NxPn8BvnSwHYEb6XdWWgoKet8gpbpQpKbR
TWhqPFU6OGePqZwghdgq1a8SVcg0pn1OOkh/V1c/QoFcF2dKQJA2TohRlKFEj4hZW2busmzgS6K7
gehPfOb1n4dK2mM+QPBRwzn/vn2AJJyltmi4U3J/ZH7rPNvQJDMZkJyuH0R6QHKi/bZovH3Jn2Tc
jV4d+mSP85epiYgOl4il5e9sCZVUbrWMkh8I/K14cvtf9hnwra5MvTh976ax0vl8clwpqJNweiCz
hTyL3l9NZPuF2ypkPdOqZEiSJmebY+ukuyeTUi6ZVxcp4qK6rr2ko02dv6dVB3BxBvgQv5delMF+
Yn0TXt7HnwkmDZXPSR6XDWWHywYfP2kI5TfUSxZ9OT+vGF81Dc7xK8ZHwRbVCvOHecMR/XY35jNI
c3XAFsSgukNxIxs+gHShkIWP746VW+IlDfu2ww8qvoJfZ7QxHaFGOqgrewKPA4cehV7ZytwGSjah
iDk0zgsbK5JnzDaEfSv6TpttJUY0BpFghBfw+Y9qnPvOVIHdSKFp5jv0UBFPwldcJgFoz5FM2Yns
lh9j3gYUV3XkbGmUQ0y0A/qHUOyf6NF6Wz3NQly0cBKt8R3aUoN59QwFmWUQvfIi0RAG19IA4Y7A
bJy9/DzrIq2tYKWeLNSc0mOw/mCRwjNOEdSCvb6JBRs5InB68k983og8mvMlt3eOIbORgWwPYkYL
q/lqzVpLp+RMfaiD1PJx7P1Df3gBQ6A7Tgbxkjvx00BKWoGcVG3u3uCRS0UxVmNSuOIP2PEoUfsd
WwFR3yVPwLokKsWJEOKVgQOxUdbX8Hf1JqYZrWT9sbmS63DMO0YRk2R9DJCLKLEJ6GAGLbQ0uj9K
O0viiD8CZL2C6r7CN7AHv+94kDgykfeijUqRGEtlmU8VBE0B1AaMKeIGjvOT1dVPqPYdsArRHbwu
/nh9xEg/pV62mESt9gwbak8MW3yj4XBf/fGBAqJhSP1Yzk6ZNIfVZ36q1L3ukLsr+uORgauaOk+y
k6o/8koVn1/6y9yc16q6o9U7qfg4ksPZu++1TnU6ylBlSFW+bdielGmJyHW1f+Es1uZywrGO2whl
7DlgDJ9l2AvDLII7g60GWYTkSnnAc+CssN12Z579tEEJ4oY6qKezZ9TXCxIrfB0R1eZb9nDDjM2g
F0Ulhyy9+B+efW0k3VJi1rkzjmIFj2waUuVPNUrdid9yg40OIVtwHsBLGwEvVJbA/FyYWC4H5vlv
0Zyplapi0mqwoYt1U67Q2VwkprD9pSTMrS/0zgolc37Ag00H8Xo+8nTKrC/V8EpIzSb0+jlMMntS
3NB8dpX8mM+T687QEY+u9NijsRBu+NDa3BL17/NsMwWCh8Xkcdg2ylEjjcOSWNPKPTq5HWjizCBw
Mg0akn4w0p0K5swQzIfUjw7TyIjZh/CVZUQ+WUoPObMV947K776hakaAOqlXJ3jOjm73VWD7jo9r
fnPG37kcWPfOU3bfMks1lnpgEV43JLA2tPe0wgNNO0ZgAF6clMmmAcaVs0xVkGuwWfxtj7r+tx0U
GSE93e8xcpulimLV++4DiffKPqhdlZSPbq4ndu3YetmFrMdMRxW6wlS+2p7oUrNHyL5fj5bwfgdh
CJnFSK3LcoRC9uWPCux6kbkxBQwPVD1+eGmpF69jcD2F9rZo6+4mMa8S1Ip7SoRdNOA6y1j6oQCy
SxkQ7ztyHKmnYZeO9J/das4euF9vnV1f3BF+pc+9IA58P4OkaPJxh5EcN27M33Uv3e7qspv+ROmN
8SZmn9Z6wVKADBWcoU9OeN2jI3UZ9BGtwFxVbdCNMz1ir54aP7oARyf/lTgcJO6EsD3QCiSQTYIQ
hdib4NWkf72YF84Zc/s1DzxdZfciu6HwsHN+sP37+snWY5/8kYJFL4F3QBkhcLq521QHGQ/qMRiA
RzWmf8b3ygNtMEtkQvxK9UX5v9/gu/MfyJISl84+LpoZTaVhUI14DReyQEZLyUeA4ZhX4GgpnPkU
LK2W4M8jgAQpW/M1om/4WuorFRGFhMaHpnNVUF18TAikVhdZUdELXNG+pTBK8dWZLz2ZMCw+eWuw
UqP5RfNu9jJQWn1tuO7gWGw10e3i94UsHxYaOcnIPUfiHsZuqUOEh67bjFyM2gLyrOx+uqCDp5MJ
Nc5zLRyHCTX/RsGvYht7g2JDOVj9KJdp48we0NYXYbU8Qbk9iUqH4q8ITnIpzy4ImPeIx1//1QVK
gyfUfaCYnpzrAgGj6gi5t5hdT9EkP+M0R2rltBaNpE91VoVRt+vyHIC6oTpHt/btQhNLuzD5CD3p
cPifAcoNhJlPChu+/BGXSoDj5/29YhZHg0512Hdh3ELz1jGex5cFqNI++trXXnk7Ec3wEbvis9rs
ij2pnGfQJDStzQOx9oS/Rv3zy4Dgkqwm7jhsIFRU6zZrJjz6Z2NsO9OXDgItBfTa7r8963QDPMkW
2STqqLtm207b+qwTd8nzOE8rTYkzHtrQEAWdki0crWUCOU2B+53cc+ZMOcIYgqmgNoGAaz+sp+tB
6nT2DiDzuIyFENTE0xEN38Bh4oY9cRWHSj0Rs6S6PjG+Eixq5SBq35uOWyCE67G1NpK0qj6hNUOF
gNpoX/X1meWW/GItRWR2Ujpk3IvMLhA7oRa087eqFRZLTuYSV1fZExs+ONm2+o1xj3EFevRcCjaQ
rPJCoRynw0UzV0rlmT5f1L1ibWeE4tWuDbsKdCXhrBUa5wz3gaSmJq4wCOXmJwQmwuNuaadvLkQT
ynVhds7zH2S6USAOnVRLEE6/BKGIjI5ahMSlPJgGp0SQAk+6YvamzPx9Paqibh6sgH/4kWDjZ+AW
plKfPgJNWA08rjvJqETjw/F0UgvxEfFdYJ33WLx7yMJHxyeyMLWN3HwhMx8b6zkYrOcmm10zPz1C
IuI4legZ7KHNPTXUyUd1OhrlRTFyfTRN2YTkClX45QlwbUZZQVEgsXItUWjmeo7gp1aXKWGnMfcD
YFA+NseQv7FvjLnlyoCffnJe1li/fFsG3FihA3krrZ2YO9gqn525ImMHiUH2etsNHQEUM8uSI+wV
dO5boD2Oh7gBtLQpkQsvffTBGuA3kc3vyEJx+X5V/bIynWOo7R/cTjDkjNiMSQuRzv/BJ6RcSMkA
rcC7sfEYL8UlypwmqN2Sf5oN3uuiuOrBmRzjOKm5GGnG/K1XsfUTR09/vY55RGhxqz/9kUbneBbw
kvjh4tA9K3Q78W/OHDk5wV8/r8AmadBFwweDQKSjTkatRHuNiC/4J9tJX/XAnQ0IhX/o2MC9cL+Y
ZLBzKbQZP9GGS4DoJiWG6P8WpBwVf6qzFfUiw+bomBOKkya2Wl0KegrS1uOQkv5i+PxPk8yJj/Po
S5+e7xRGD/kBrKhy/MhxkAdEF5Q0Bxv34y3P4CA2S5EfJFXh4OMUuzAh+usJ/uc2pz5HeQb/7JV4
qZxFkw4VeXXj/jQqQLEKwNS1jcuNK7FFEc2PbsWF34KR7x6cKdqOtD34yVY9YzG9eO9yniLxmkwd
FUTVYDi0s0TITuQAuZ3lBmWInNJaim7T7q2hkm/3ZFE4GGqvapBBXzVuPZa8+fLB818ZRaKSn6ze
18uprqphTi3iyt6Ml79tcYlYW+NLMdZe29vuJSLNNbX5b+u50srKCWA54XNeXhGeG1DP+5BZFZ/C
GzYCdDW1USm96bJlfDgZYM1or4DmcgCt38kQVmllG2z2MzbLLwQDUC/WFGrsCRYrOb5E9wzGb+F2
cOwj0qweomSX+mRft0gMZTstbMVEh8JslprCj8o1jZYIZHzIiVWgUrd7BkHqInP5lYb2O5jOvh/B
tRHLJgUiQ/Wpti720SphJ9kW93fudCki+bpUtuBls6LXdqCmWzArTB3LiAZjljRovUuoli84EV35
IOjiYYVjJOBt4auIC1ezOu5mqAlxAA5mimEDqWovkIz08qC6ga/W6L1F5L9U43V77/Jt18grh91l
Nwe/l3n6xf6gz80nlPQzDO9aFCPfyU3vdJ+WOkRS4UZD22Tzl9sE1aIjc6yQnBXZvhize53ovhEM
6u7Orzv4iFiw+gh82iLC2BV7vf5mcmYef+QLx4RXlv6q69RLXaaXn90sJiIfFMrJepFjz5ZdQ7DF
UDuyn+6OLn85uIB6ZYH4296+apTuoLCUBJ0whFXCaJX3jAxsy56OtNHxvsTf7TN38ZP88HBiPzwD
w2FYD5P0LSZsqcui3qeGYXkla00FjDBw5Ip4AxVZXsWJjQccYXi4F/tfgPANWLmlrdCqkqvgyOWO
kj4aMNB/4gDg7eBFSmVH2NlkimgbvA76hbsgevVs9TOteUUOQq6uKMhwLvWnIvKXvADPpEuUQDpk
0h8ELwfSA3SdUiEEn4t7SeFojPibiwZ5NbgpNHV3aXqcp70bjOCqfXX/8AmvGtlgLTIPsX+n0ksn
jHcYLTS4U6epORC8ItOb81iDGDlPt3zaNf9nmgNwOCmk/5ckkwjAzBo/F2vkrHQ4PDuFulB0wTkO
p2wHtKkJcYS0/ZNpdNKHAnl8gSHB44epzd0Db6jYQRtxVvE55e9YTN+P+lJLc5SMv2M9rAH4BA0E
Y6KAVtX70w5RekVWsUL9rqo8u8wej8sby3mcY3/aEdFbJSaji8NSTukB6GGIe1fpxThTtzN4BjEa
7an3gV3P2kdfdCYcwvQVZ3MrspZKqz5EI6UNJi2vFTsBuaVclgggJBY8TfQUy9veP5oFf5hyrvQr
zpEb9OAydrcVkcBB3i2dBbvhHwH+ZtYg0bfzUXvViJUhJwqDPHo9107DJ+JwoC09OFIyJG9XBcyj
KafVut8uKRJ0nhkg8VkgOar/n0ZxYGV77zwz+EbGkRNoxuB/mlFP0qoPGyKCCExlq8o9fBXmBsk4
n3RnH8lEG44Z7qJ+qnGlNEt0fp43ukpLxTpLlG/Pf3YLnufrDqqI/uhPEm1ZaxQWN7G3YlxTjbcU
IEKCDQ8T+PDhoM5DPUIhmZJNmxKE+k/x9xVidvgXw+/U0OZfDsEDdY50Hkvt2pOgW3RCfHgsp8fg
XPHiHPK+GQ9Y9Y0ZCsCavHlWWpTdZC70SCqUiDJ7/ZfVDx6KznTeq27PWnuI3vkPA/BH83v5Ev8V
DU4zdqnIzfcTXxHbdPpQMJVkHHUdQFNgVhJZkgPvymNRRAa8QsCn1uJAhzq/r6YFN2lPmQctmTdK
SDWsXOab7CgiJEg0BqzARC1gHp9yQFrwVBR2MuSxxYnjNsTe8R4XIV3qoMwnIVJEV24ajSkuyeYo
joRXDhiewFfUvC7mWlcueRa3XRWhQq2INd1dIbknIapUo9YGmzKm3nc9dYhJMoJt5d2xdBMIYAK2
13EtLZLb/cql98NEde654vkSz+2r12hAmpn9doaFCX2NwJQ7zulmhjLfEz88Ndy8/Y6B5c310054
Q8kby2NpHPIq+Zk/WxV5NdvD63A/ABRpxfmOkJ8Gg83hNh510tmp+aPaPReFF3qe6r7tVJfg5y3q
bJApCG8K8Tg9f+hQQ0R/ATnA4fF9skDTNoYZbgPRk3E6jgtBOGk0S2uM7lZfPunnw0LxPmiZB7+Y
eOzfw1QP60t/6Xysxq51gAk5zNCQovkB8bXDw0YhAxvsc70k8ejWfyQVCVyAnG5BDss6lE1elhED
PilkydQBg2WumJpG29Q5c+dVNtq33XOQByWUL52rF9RWZQqR4IJnyqk5D5FgGd5rgQu5WlP6Iq0r
CyquYDatRkLpQ0lp2CJGkcF8nTf/cWvT1nWIWoT9p6/zqKMfzEJJ2/yFmUO4sh4Gdrxedt3P1RQt
Y/aQIa7p2U78DRgiLGoCj97g0Bjm3bidkL2Tbxl75UqcYTEVs5EwT9PeSCP84Ce3fKx5zIR8rmHN
XeE/IAiMQHPiueGiOumxPuj8tF9auhKPJz2SBjF1o6zowQv9yXqZ3un7LaxUn0YysVm20wNgvE3R
DL9F3KAYwOyUQD4CxKGN8T66jOYuKsUcMr6qiwsD2x6BsUTUsb9jrXUvx/NL8727SYmZaCu/98Yv
fIVjhkxn3ekWtGUciUgq2KfXs/I4v29S36E325hw3tm/9HBRG2ib/WBgfHF26LMGM8ojQVrTE+mn
Ew43uq6hfO+h8OI/e+X83sIPFjcs9PjSGyytxVJ1B1bH8UJj3nwunD5xrejbyDymEbxn6bOW7WR8
BhgoMDHHbJrcaJ3TeOOY7+ZCQPdOAtpRaxZjTHEd6g97Pl1GcWFIyCcu7a9ZRELFq5GHPIMv2Idj
hUUdoPXruppbG59lySo0NQ9XJGTaHlZlYZ7SPYfbplXbseGAxJPGvPrKdq4WeSXG7q3JAo7661d4
s/1p2aiyM1T0Mc2V7MHWkg48nxHrA5Hns5HUY9e8q1r7aa/QG3NLI77rYIqQk0i1br+kGbc+/qn3
LnfelBbw3rxNVVnxwnIxdS0xqsbbI/OTTKyw2K3XUG7BCxnsDGCr8IHmZJt+cCavORFclhw13aG/
A3vnytxV7gv2yE2wvdQzM/EUhNStbh8QSIA++BloAck+alsiiMTpUlmdWv1/hnTV93MyiAFh3zRZ
gl4ZWQsTNJD2fqYUaynDh2OaN5TVOOyKe6KXQ1DxF/yR9DPWKP7k4AmTxTrI1a2gNRmCncWXT/NI
RykWqlSbWbt22yjEtoXRmFQtnWekpgRcY8gp+38uvz7H1AIXsFCBkcJihSKaIQZ0zj1ad8Q+NOYE
D4Z8qj2jafdKd5zTE/mYYmX1HyEkNE0tNZVAY2T3xehf22on8jQ3itHizbx147mgTjA8F6In0sdT
Xmla15AtAL8CRPaPMpnrn/jYe1Kgth5VTmKXAgcaqvwWlNSt0KeB1x1itKJCKu49EF0mVxy0qMM9
SHqgzMoMSLhLsnKjiZsH19K+CqC88AwsxIIep3Iwp84NmBgnilIOqpcbB1RU3W9LHgzHHsOv8P+M
7urz+PPDVgelyM2DgXs54ytJd6Ef11N7HDsR2i3MLgYeBhidRLIKzEK1AaTYGR84wczH8Q8EOIc6
6iyrQ++VycHyOT3v0djw2mLC4KTTIqtYmKcK1dOWPWoBhIuzxv4SgWIh+LWJ41dx8/qRmBdrRbXX
iCk+6yUN6WTAtXoMK09PktUhI/1t4NnCU+fGAnQYbyjP+KBCS+dOQoJ0rRav7zRK8LTgy7r3RIbg
alg3ggJNBb01mozNJs9tkDC9WGr+Fj/hPhPu1rxVctZpYgBLyVrYVDAfNZgi3xWoh8yU3LyzdY6g
BPmZs2Ngry90u9gyWPT1KpGoPC0RpnueF20J/iYpcF1kZar7RhjDm01y8LGm9/mc9I8cvZGofdJU
VSgQi7CNnSBTXiq0pynkJ6fVcFVDEJCsn/WfpEzIs1LXloqyMzRt6U56cmfovPM7yRy7wjxDFG3t
xEytM0zEWZZrA+TkHo/PK5eyT3/7HeXmyJvgyUTAJZrzPrN2MKjvfzLaizGeAse7CYzpNf82CMj8
fI4+4AjnIlFxDn2rXIbDO6anr4FaxhEVwzjXQBEePBw4uCjQRWUPn9k4KRqElCNFkipOWVcSyW5b
dX5g26V5GAqF2TjMcbRB9DqjVLaIJ0QfOPoRDvS1qpw9UTJ+1YzECYCf47A67jr5JoMk2Ntlqw8L
qW1bnrfqBI+uYuAAIuyrK8x9UwJtM23o61jN/JCYALH8fPobpWLuvUZkPOYWXz+bZnISUSGkaeGo
Hmr3zlqcPRGNvK8NomIOqVN2m9k+kfkpTNU1Jxr+QEfZlkBAzdU6h6jldOgksKTDjdlq911omaii
PpipjJvxqaEmveJwKm2whiHlnCR1H/+aZ/UmmM1g1e/Z1TkjWUIvxXYcqEGc4tqkyTTh6wpNNsaO
7xBdp701f1wiywl1GVj/D+Am50zOQFaVOYC7/BWibijyA/o3hmoeANwLxFHpfSFR8nFi1Bu4lknz
HDOZG7Cc6MFQooT56yXvmByx/hcKuHC9nCSlvUXNfUjioGedDZldPEmilAeVtNsU6u5spF2HbCED
mdUBHlQTb63GH0raFgOnyV0VDwzluD4Kpol2xV+tQ0pEKMqiu8fb9TQZXcpqzgba7rSup020SWKo
u9NIL510/pg7khyn1dCs2DpQkyx/rtpd/LnTJs1S3YaBHWwxPhbvvjUtCuDrBzRxHis5Bf19k4Jk
xTHA8yT1R9z97yn5eLYTrScqRXwNTIxfols+5osl2FovUa26519W/Ki0Yo5IyEcfT3KBuL/7rqp1
8z3Ywl5joCoQXxGTD+DFYSpOOzy+XzcQRLcC1U6qGcEj4D+HV+iJkYqhkIHXZ7uEbiccgqMLGw7K
oYySVuIIXYC3pBka4GDjhejcL1h9xNr+GDI9Z+iLJSqzYPqJpqMid0RMVpM11iQh8kugS1NcMpmy
2/upjuvAlBaLXZPVuwJcLeZQ/PWSn7AdeI6trBg8lLW8AJ9pWmSzZw5r/OhY4qLy5nMzpCg1iyKu
XJTfNM8ObNnPjrCvjRDz9/xxnNJ60ToDK6EwBi4O7fWNtyJbwUnEqj39CNut6LX7YjtAJ+vasSSJ
iacE8269NWX1EWGTuyxSrVTq1FKP413RW9s9Q+cJCTYMffyZBCy911eLcQORiVvPrgBjpyJLG3rY
59RVX9JUzG69N+X+8QoWmMv7Ox0vuBC98KHHK9VQQYksFecnmUACKlsSeRC3U+X4otzo8faCyfk5
bnN8SkszZGHQoYaQciIsWz+s8E8Mc9bnneMfh4EddCtZlzVJXp+bk+xapk+Uc7khEghw7PA3cYyn
ZX/v+9xqhnQikhWlm3f/nlD6aiDP38Jv1eB+fgLj4ysvRyCIFVerhhDz2937JRAvE7Y9ecBnCLsw
s24lp4oMXfERRboKRkGv7ga5n70P0Je22J6oPt9/JNDwAWrwtQWxRAcnB1HqthlQPgxIbmkL4I/Q
CVQIA8/i6zdXqGzZ+ioLQjRLYTmN2WTnWA6C2BnCR5RzLQTNAPRf3OZWoUbgSGc8ISjYiDgfeoW4
SZGM13QgnjqOHQcFUmIF+ibW0vMGpytTpvwQjw3UGkths7Q+6P1iTUokiaDesfU/A3F+5dUdBP1z
FuYYbNsfZwaBvHEzf6LKrkiGVmIHem1KYIVU1Due0cWjflnUd2W9wL1CPoABbFTe9mMycRYdYWEI
gQADya59vIK8loDIGvaMp3AoGodGGUQ88xWQ0jH0Er7hYPfvfwNZltt/JJCg0zA2kClf56aL9AyL
1XWcvpqiKW9iQpG1fXzG8QJvsDiLHIEFjbuJhMsMFW7EutbmhR2BFKu9c4psL6SCkaS/2EYhQH8v
Gf1D5KswugiSUOCNIBNZzrRP4+J1UGP2jaHHIsjXCR7CzTyWhk70Y2uTtD/jJ5I0gcqORpRnzYyE
+O9XYgk/uR9XeOIaxigWFZndFOqKa8in0nOil3na2IYpF1pToi6+cQn6ZlD+RsXLs4hIGPzsLcFI
wJbNyFSlBllmbLqf5IYs9vVbjrep+/eS83bm3ok2NY+BaR+bSOv7cg9SkAW6URXLZUg8sBUGsRfl
Sn6JNOHPCsySAbdXWl8+G8O00mDmfT4pfUoGSb2PakoP5Ayi0RzF68/21/Wk8IpnRPY5Cucdjs97
vEHGWuWEx1E0XE9R4oFUd3H68+UBtiOaq0KzUSm3Fu1zfbz12C7BPK7XUR7R+Vu6mIr8gdwxJzWA
nw8wk6/3aK9NpBOGrpGHl11SqmIzeDkxFHAq3uWuY8qeg/Ht25+AyFhm6bZpe2E4iYLLKw4iBDCY
ccmVfoK7s4CFGgLfr2LlrVjwGhObMd0PawSTAelXAfB70elwvsnjqQGS3rLDpHdBAe67awKXbqC/
sPDB5cITIhvkT1EMVorLr8+IHQSjDCbFpcB9U2Cjccfr/GZcHwU6PNYvSns4tEu7kAqYch7Uu2Ch
J0JjLvjuQfgbw7V2KPG2x0pItdS3Or6EquXmOzRHTBz5ib+/Zmzi0VovUek9kaAxzTxR9oGYlqv5
IrVrYd4MDlJB26wQaTgPqlcLBER9hRPblqnPh6pvgFqPXwB5Bvi7L0tsY5jac02fTnvV+NWuEv6W
w3370uN4fOX+wYCT7pV5kbRJqGFk11ITdA6Su0r7eBb1JAyFPPDCWE0dSUDHheudV6A8UvyDwSte
pe5Dg7ra4YOb2xY8stpET/9L6qmzp9+faYjHh6DkHdr/xCD7AZ9hOxd83u8URFb+ghJwnSi/21fx
jz+MWjH1xr+hWdjEE4B5dZf2KsFbmHGFxidECW1B1zuOnaOTZDelwrDUFMx9gYCNxWjsxZ/oEGLR
A8I6koyzSP528O1qAR4uIuxPq8xTrhSSLIIMcIYlqMF8yLheu/LOI4eiQHd/iuFSXc0bh75l3Qwh
3uj9UIpM/v8w+DyEUTKhzu/2P2E7gf4Em++UjaQxeVsRkypJsxWhip7kSEkUZGh5fmnJu4vfL0RY
UY/3snoLZpuIvYdj0zvX5KwyQAUHq0avU1Nxgtsjka4sStgLx0SdU39Z5XsFZeSAT6MLj/MrmqhB
zJnQNrHtPDqJboglLOdHNXktP8ao0qIcF+KGINHc8aOLxpfAyQRALgfHkAY8mhdPS+ecyItAm3iV
ZZn02WEeCqmbQDKbSAK3Q0VDQUqIGu3uiJw6EeTDK4bhmJbhc7Y7Yvtbv01TaB/75fOpXz7CxFEX
MbruqD45HSLsTZdKV2RO7vx02r7W5GGeGA8mECtloZqlsQz8233PbaO/3My77lbUBcb1hpbGJgeQ
6TEHf+dfIL+eCp4OZRr4BFfh7+tts/8vqwc1u96kE+RwZuSOz2RPNmGgzlXxuWVso6Ivwz2y1nPK
oyfYFPdAeKX1nC3acFsJqOK6Ibyf9Q4hBBsK0Ug3QEInOdMp3USHfpFFot9kgOr/v756wlUofzXr
FXs+voNKjoase7FM8bPg/fSyxeaJECzrg9pEonxoK01m3OykmX4hyZbkoipw1CBJ1kgG/gSTRtDa
zjuhexJ97J2Uve71o2ns1nWwsK4d3678GIUlK9xKEMkAxS+okXH6GEpMra7nnhReFoI+QcLogDPt
Pm6WR36v++RCecSBUwVh0w9zJNe82K5u3RDiDVU3hbf42wTnoY9dhM7tQP/CMdUp8aDvl+tOEW/I
MSEYDV30k/NUfm3woByL83iGCbn9XrO10dn7xLQJTc7Q3sxWkWRq61WGmEhrBSXm4kRmAZL/VOSe
Legsril48DarkkW5MdyOAOdtUDPWXRh5sAx/AS3TFrZ2eRNsNRwnllHfdGvJ8YxLZJpkX51hh8xa
kLsT7WXQzqZ6N9FRQkwf+ZS3pFgntspbCZWUrtCw0A/VumpnR/prhqHoq/KGfejTy83NuJWASrUP
l3HbaFcoBptg3j3F7mncXCjgObw5U1YNv3sfc/nI6rFVRSQyReayWfZZZkMgACRbdOvqibDQpUv3
FF9mL77ZimUC04j7ERfqq4zD21FcbAt+rViMTXRkr0s08Nfgg5WP1bls5v7qYot6aRUTzoy5mRwY
dX05AJ1YOy5NmMK5aFjL1i+D9zM+928fE0ds+K+MVaYYPuEEif12YbGPzDkuF1s31hr3Inwr+Iq8
y6iWTbSYF0jXZPAFJ8ZmXyNQfKX60CxGw6HRhyj9Bz2DA+d5X8jHs61qDXyiRZBAk/om8ZP1/llu
wRE+KAsLMLGhg/+CucANwyIDT5ce0zPpIE16bNvd8JGEMJlTKHBHbgDnVv7S4vlMWFe8O7xLY6hV
8e4tYlFHOGKMHHq9i0Y/l+8kqLEqxlooV765pbVTYQCQNQ+op/bBoH23AhISTi6BPKYkK6rh2fLQ
hO5O5f5lR8jsIger4LlxiQf14qg62Secgz6c5mxzT1lRu8gnG4CyjO5dWZd/Bu6BjHrcc73GElLt
khBm+I1bLdftYYp3jaBunfWAw7WE+yQNOFPFKcHEWsz4X3BCeSl8IQCz6EtFg1qfnwZbKXhgv2zO
yg3thAa1U6J1zkl/xv0sJF73z5qNXqwvLnAO1iEMTB8e1XT1sGKhRTj8KKcCAVOf0rUEcpcvYNLc
H4+8r4Dh1cukBqo93EO1z1FPcvpxmUi8FiSdU7/jSihuSpEn4ZoiVmUSLmxzG0TtFHolSByNRaHc
uWS7EnLXAGpcXtDX5Wiwldifi7DcbXlPGxJj9lx1zxhj7vKPDhq9IuO6eibiPArjOKBbbbk3LhAI
0BRECBF7r7ZAfQ0hKyUCYyARG89zNfNH27WuEjfQsD5eECpFsm4cHEf412crkg7+hx6G6MAEc6Ev
tx9FhjN3f5VLqZZ89rmQ1xZkG9DeH4+YHKMNE3HPNOVsfJIv0WcbnNIUn5HjObiKHud3IM1ExRXB
uWsnV8WoA+VDa9STTXKz1HuPNvXoscmZFEZYMza6h1JGRNh1A1HOOwgxzBo14eoCxxhN8cS4F6s0
f5gmAhSR90o6ox2Ka2yw/u0iFAwvdGA49iavw08twkPL3KnNJIMlG2vvSSZwCEbM+9Jafco/caRh
YdydId4e8B0f0IQJ8GWWWJw0+u64JifT0+ln2+NlyLs5LnbVrzKWrlodqA+bSDfDqqSe5xLbFSxr
8+HTADXXdue0faWEKpGzetOVnmltxfx6+DuCjp4R+j90o4yakLASZLdWAupYIziM9scaGjxv8Uk0
twLuy5cEnnA7jToyhSMSxtRygtZTmgkfkfCK7N3+iDvcA1UcGa6MNSO8eaxjEMZrSQ1eEXbGANLI
wWNf+AyBOVkh4040Baga5zFoJCGaNqMVtiay4RLNTPW0VfzoTJIEYfjq0BMcOpbJplHs1YsiFbfF
R7GlNaPhG9tEvLiU0DzI9NVR40u0YWFUP0H1EQvfbxRjEypUrZ6k5E55PqvRb13eUI5js94COrNi
4LtPEBuPXk5iaYnhHbnbHA2vU6tgRnNSswzyEdqSsa2RRC5LJzXM83QmlGgRV+/LtigAK7D+K9v4
FmIXaqkQi8kLCPxX24KCjZDSTXNujYJaTPJNRYAlW4j4Ce701fXEtjykt/K+WYLbESZpuYLjUCDW
sK1spTgCkS8gzasLSG9xh5TgN0JZwhqitKr8t4iU0RqhFuEeyh49RBTiNQQO9zlqxUGhGOMrYv5N
LOvRxKIpySCym4YPCVPzoeBKSBg0bKsQsRIXAWkm1DxEzfXqBtiTUMhTsZGar2+eZlk/LjmT8C4z
0qBz6tm/6BtisNo1xwySn/P150ZMlPqsBn0HntGfpR8rAN53oPjeFMwfCBJrKbu6o3j6IPu0bOr6
pTSBMlJs6H0u8QPrK8y2DPt3DcmP1gX7qvw+fDYcUSjsIEwdIYwSs+6jLRq1X8tWJYs2xsM+EPKw
eSRXeeuDSnI+71osKPcLkNV9tDemPUQ131qwMDzMq1wMN1kpnBd1Esq978V1/XF61X4xCTWmxnnf
OjWpdxk1j27Mb42q2/ZRRf+O1eZQrn6kcXIFyWCxuwqQG/AhNGaB18EHXAcskHAV5cuiCWI/kbru
kc3jy/KbkHHUHASAV3/MtLpysPc+E2gibQQ0JNjsAHQgHqi1Da3oqIr3mmI7EJrbmhYAGbMRdc1u
Ln6wUeCCuxqdk+1f+bzhNXrrzupxPHDixTTI+ayL8hjdNcJxTPU81FZNL606bchEcxVoi5SVzvEt
LMZW8sMOxHdn7sXUH2nKVgw0Js41hcsW4xgoHCueiC4FAE+vJRdqh1j2zZ4B++vgW9hPX+p8vuqf
8AHJG66wp+miagpfvMZGke8uyR5AmxZP3wK41cwrNqGE56IO1jGvgLMmkszai5RvTUCmS5XcWYcX
hCL/NsGqdx8gAytRATJ+rj64TWZw6FPwABeZHH5x3b59QzSVxtwkerwmVqIKp2mX50iSgRPn5SLj
TTJQlvgGSA0olmUZFhQ01gIJeSY7SM+fwW65LoZJ4zexu+fd9SFKDjCgHOPEWOr+gSVZu8bxeK1I
+JXZO1+IioqLv0fSROOTXRZHpN/xoGnqSGtGF22hDtBNrjbWm/qSAD08XVb8ZsY4KF0A1KqE0TbK
mjIpLnUuIIwm1M2Bn2z2sohwSzjfwzwvP6EjtIG1zexoL5Apy5wSLF/XpqbhQC2AJEmUqyhCMAzp
B7on5mhQnvhUzsFGn5a4w9X8JGw3JKmaRrcCuZxxr65cCC7OFXLtcB5p7q7ecg+/O3jGkRMrqCC3
rZSvYpth/mVJaegJjX6a8TD7aGMsbUHQjJrJuvM5mRe/7QGxhxLPC69huidxo7R5xL+F+q7wl3wB
E0mzxMNIILC+j3PXNKBvye3rCy8DYyh+2renA5rOrLc388/iS3WdtPTK3XldBblY71YGYvjfhNdR
c2KkDmIKnW7hqs0wQbsYUrGjn2dmu1nc7N3VpV4+F2QEEhpUh8GWBlJd+S8e4WESED/f7aak0BQj
7oMsR6nArfjSWu9jWxLyoOVV5g1+fteHpeXKud2LLZzObN6Wr+UfpWwn+yvS54LPQzoT/2n+dIxu
rvv1PerlIO4qJaRlYGg04jrrVr7XxzJi6oANrYkZESFUQ+4CQC6TXF1V5ffgHZZRt6FYf5eU/bRE
mXxWRIgP5lllLxBX75+1PQJFl7QEtPWC+11vzfRhThD2JORQhi2niJ0QhUwbACMP2Lt81uR8Q6EK
GCHTiWBztNV36lHknmkTCfnqyM+V+McjqIOB80HRKubHV6aBwToxEuw591vOAXcUyXa/HQDIO5M/
fWJicC/dolmo5f3WVwtE41dYRFz+V+J2EMcu6I0D7Il2P6g+pWlEaCSX0KeNr6NMpEsdkTzeg/zD
yUsa2nxbsM41u0MH2IsRsN2bYymLLY58CI/VDNwpQdllAdqeXdoVEY2K+p6/2Y+ozvbGnych6yXX
6nMmPUHc2XjtcDexx2Q60kbOeA0P5yMpK5oSmSIaR865unjJIX1Tkx/zjNkNpywAZMsOEfrmd1ES
T1O1sYDdp4TQ3+lVjG9QNX6sljYeXsuvXlU+QceXZdGawD+R7h9sbYXkb/v/7hdiiKNcimVU73MA
w04XmHeRPem/NSEqgZCt1jBBoXtmaLx3/qLwUzjzEqTfgEsBp9G7p2aXVb3QdZVPyCB8LznDjRQp
FrT66NIbg9PBLm0sn2EIsbDJNckhAAR77tIB4huO2Oth8OTAYFzwNc1s7zeHH7Zrh/vY8DtmD5r6
j30vIx1HFOtxrtkxPe2Z8/BDpTuRSOMzt0qKT30RiQWJnEWVhb4cc/C1tH0GGXibow1TPm5JYk+W
L9EZnJR/j8IqhdkxNXEyRrGzAYLKzVRdKhheHO1Yd/T8Ojla4cI7rTytSbDfF7xt4QIw851j5tk5
0pWkOWY8fIFdsz0TVkD6zINaEhGMLjy+fi55hypFjX5gIiEvK+tobkuz5O6+K3B9Rf1JX4Mz/9Os
uoHSVEiySEQefH6KynjPvdSmp0z62wmOWDvELIKfa3L4lo5IKwr/1M7P4GwzN0bUZvaD+g/U/alA
EWbGUnPKkBx/gcUow3IaVZyaXjxHfY/C8TINj1OUAEU+cSpCEcu1mgJY+Kzch52PTtk1geR8hd6B
/erKR9E9jLXnND/K+zncYZTLRrHCOCAnPISc0z8GUF0PWdH+RLhaLyUUXuIZjR/ipzcpuhOTiggi
YxllEd5fb9f4BQzpVxC3aJDOJCkjd1j08k9PKerFiYk5wGKGfpSBoU0rDy56QrIJTcitUHUK7uNz
pXn8futp1KgGNmJSM1Prgi29j4pcav3fDaTICpps7V5GRywYuXoUa1xLN7fA1BTrBPVxNdU3D2hy
HBuhCNMbCHReUzlNTBm6Ldj7DDfpF3g8M1UrnWazo6ajzDY2LH0vn7ula1dbvwYJWGF8y8sS24OT
6duLTa+lw5S/jWuDW0eY5efradvPO94ecIyaQb0aD4OQHZ1AqcgFuXMyx5dPi2Hy7Oscq1EtF3D8
X71/nSBRib3hRKozU6mbvSoIzgVg8zZraa80UFofzRuEpxffJMVOZ3hSmjn7CkDOVr0cY1Hj60IY
WtppmNMHqUjAPj6ZT0m0AxqFQ/QjGBeJyKavV1/AkNvegvPJINLa/bu8iXOiutmemUkkP/GJa6ao
dnn74hu3oOym99X98oICyyjEYjdpSCLczp9eFctKqLFDgq9xloVckQaTQXiheY/MRJ5G+OWrVI2C
Y10jm3ILnhu5nSMpDWdWKg1IAo4vbOCRCgQRf/f6dJr6lVInoU+DiL5oOVveg6rft5n9VMqbggNy
qUjLFgBsWxml828D7mpXx9nmuQtbFXCTGTyrrYFAbL8EbKH8xPB4nlkhGrBGzcZoZjsTS/tls0Su
sKkrfZShb5eq1aH6D5PbKOGxMLAzcLZlJKg/oK3ArQcLfs2nDXbDmADilkY2Mr5dmOyqUaiJAc8l
CHNMfGESkr29R3Yqt8Mp9iEq93MpzKAjpNEPKAZ7hfSTCFkDcKOrUVO1xJ3jGLWbl3KWuT+Olyca
eMRKZKIjqDr2VrH8QSZ/mCQmqD/evNmoR3Rwixx+PU5E8M9WV3WiyVzfVH2pJ7YCIIdHPoP4r4uX
gRIh/I9t/MhfeYMJb20FpvipfhA5vXd9yqtaxBkzdEtKSfyJzq2cqrLmPhk/OERFYCDBHGNDDSP3
3dI7b+4w5wxO6E92d/DdYn8kuGV8xKZQwQ6f62Ovjuxi8mhpq3Kbb97H2GdoeynqNvpydFRa/RGu
b8u98QaNGH9VaXgjzaAOoGvOZ0VcnBFzgVsU9COtv48B3u1IRKEAOaqqrBCv6ui0ddWiFW4IJuhe
NH7puD1cYJJD65DPjjMMEa2u4wtqyKX5hamZ3WBGyiqSZulWPDhnTDJ6454nchA7hB/9Afq3dhqX
flia/Gm7UhyHMKBpDWxu5KjFz1Bumy0oseziRihtwA4WN5A3Z7bVSeNG5UwcjTIsbGuGW4LMTxkY
pxL82nsbaHvNHOLkeqzTCOqudlNScrO8ysbY3uRAHVxjs5u4lzNk2/iK12vTeDdbQGjYOWOvsXhl
ISVQ3EU/ElY0lHgOGfvAIuDJlBIFVGfbgghLtSLZB6C8W2JISuWfpAxW/4OZyY9M1YHiITSKTIe9
285chhHHxb65EDw9OZBJdQ2eUcVzxjA4Xunh8vBl3wpEgxvgy5F3fwyR/dYEP1U1SgTG+1LMV4TV
6LYCI6YjlOGm1HVZcvigTD+Ksfcgr+sSQcS9cyo5hoxF0FRpXV2WufIDYjrEYSlDm5R+kmAeB6Dt
nPx+hM+YnMYz3lmHtNu7/tEyx4zuYys2lMj1bKoSAFpNqUaPDJ53RDaWNWnJRlFDH+h5gIv8byth
ROBJA1ae+bzl/2Pf6oz3QE0bmHnhjkYCLLNrOs5yHRjSZgC59Y3RhW8QdrEH9jXYZamSlFRav3wr
7/ksyDOXxMpJ8dO3Kw1/ybXQsm9k2JsLOSdHC1GdMOSGuZAV+3XmPCUCxLquhz3gNu72i6a2sLqU
Ex22Oic7/HGt/m5xj7IgXduJ+xoUMPanNJ68XJ87PbAl0yJp4LiccQMWUz1YUh6XYCYIGT/8c4dr
uNzIYLoMAC2ZayV9Dw6ZgJGR8Pm5vJQSBi8nYMdUzwwkxGcka1Sekltov85TFboVAPQ49TLmD0YB
gst7nUWamWgSwduzt1EruWqQZSAYnzZ57RZw6OCz/oryo0hWBXW9hRB3MRELAvSUjyUoT+tUJyJC
gI+CSp8HH6L11VmdHiTL6s6wZxFZ9nzII4mQpddsykMKWYeC3FSPiSHz6qXzAdWv27KM7n+kuVBG
T6y9iGgcZo3h1sS7E8H2eODNvq4wby9niKbxM9p0AwFBXBCcQ2i5LNPgGNubRxKsBvpJiq+KDRw+
AnJxCbl34+4mfv5NhPYfetPZNwtDWNrbQDEOFcM90C/VNQ9Vi/ix8chLnOzNTB7NSnU6MqoDkJyy
G2HAxRjpRBHmSkP+yAsHRxVQTHvm6R56HL6D1XD8TZ+4iVzAPjXUMZaRfmLnvwbsgLgbpClHarLi
cBy9z9QdXH4Nlx94vH1u4mPmeD0lDDy9x7XHuNhxUgY4HAaSp4vaaHQNYI1jrw64uQNHAV6giD3v
3sl+s47PeWknwouqq6Wzf86SlgMnNwP9EKU1cCKqiSvA1/WHoq1s4om78pCTwgZG36Gaq+fydtFg
6YszE1oWLNxNBbTXOf/wXlVZthn4Mk2ep4HubBJ0qnffKuZMQxgS+GKEbutt9bxixaMudS7w+6MA
9YS0Vq/1mTwkL01zW3dA3ik6vMPxfPS3xHp/qhgygG7mgEvcaIxXAHZWC8Ddi26pSn9JtbRYaH+8
kFKuUD5CPZHfmACjgQSyEorTGM1JPwYPzJRWpYY0+AJZy5Swa7WoS3xE1ls6Vt36D9drTGbdo8cN
gS3BGtExnQZKsB3gNo7vSbsa+x0k1yG52UIZeXy/Xzs8YpIjWSyRaAiQooSP5snyRRhzBwicUyDS
9prmF+SjPrgj7MQxGY9qxL5VeRMAz9w0CTwDhW3FnQG48fDg12Uch5tWZ3IMNXb4qxqrDYwHLxVe
G3T6Jva/aiNNTZQQV3ufPA1Eye/yMUZ5WeDpIOnPLfhTwd3FgrR+klpryqcjYeDBeT34YBWsL9ra
fLo67zGK7Z7xW5zKs+kg1Hm3tXLJ/K2IHl2V2xgujd/gRy6h3514fjb6Kx0J8WfrEuAy9Ia9HroP
U3ovHaHAosmlAP6EWo6gdR4Ms6+M0+7bUjggw3RX3WqhWyALQO6vQqvROmk42nvFD5Yr7vchq8x9
SmMrKnwzPV3tBjg21BwsGspC6jFPXvIK8TEU5HbUaiKS1SLst2hSmniRzj8CMOdMtSXRQjW+HUZ1
dPHkVCEozoqTavo+orC04uPUGKglkwx0K0kWt6LR/7d7p7cghCwgjlhV5clKi+WdNknIbBJrkQBH
WpXNDDuA3IdJlpeLjRcigXcWU4ly0FtJJj5JcgNFdf2Fegkzq9zeh87drz4d6JCztxmUFlRk4PWG
IrnFLRUTlrBJI2EQsoHh55ZkHKeh77/p+DKdRmNkT1CKbgxkLHOOTx82Nmo052ziqUTZlmU6F8uL
BTMT6u5H75YoFl9eNyCYGDA2pZ3rSfQmTCbKh6gyc9GZB/e/QGVRG+uzYl6T09S6u7Odf+bDOuqG
X1oPQLIH+CCocyWbHog9K+qHqD2GZA4jTxXyewWy5D/hyFpeGHFbT4oBSptsTXIDLcjjE8Ge51Bs
GhSiembpEJEb+1SzsPECS0hDD4nCMZuevwlk2I2+au1TD+41BEdiIlkta2ga4Iry5oD7yUPgKU4e
pDcT0PkOduBzBmrETAnsJjeOus9oTsgxv+YOCmBSZtmCNMCnP3V/RX8hmkBinJbgNB7VByYFo5zh
W8gZ90LbPO4q/mKIjaLGUWvKs89tC+wa4UvN5KNNQrlodWTojvtv9c/MY0qw7g3sM38qan4hJupG
MO41Uzf1I8BlOWcOf16YeQRJWTaFhN8c/3T50fsRsHLcmjUZIZ8lD1ys6igGo0A6SaWuS6mFJ0M2
3AgHJ9cokfd0lPtenlHFUCid1IKe33uOOyoGmh2wme8qmM95zzIO8nIDrCsMxkK9zMNaLN4E01S6
3SGFVp0PNWuWTHkBZru7ugZ+i8AFGpdYaHcgENdM3XAsDWnL51wsP4dfPNMermXOJ8HhMeGiqfMh
n8FLbnI8PKEOdFR2audBU9LVm+gonagifN9psipbkBCIfrwQRuTqHG6PKipViHUT9PGmtRAUZs0z
WIscTHZLRYABpfwWIygB6qv7d0UjWwlH2eUrJ4sXv7t+B3xlJ2U3oPetZChZwB/Y1CO8K168pW0I
SryqPwON/YzJgWkVJcxGVR3MuDQn9DA6fVLtRgX/NF7FAZMXDmhECweH0yOsEdnK9Q/cilXAqSa4
yFsj4yMzZJAkhUuhZn6njQWShUJl7J9IgeB72eiYntgDus11mX7KdaASW2i4Kh9Pl2yEJqm8SgHn
V+HVCqbzYCR4vsuaIpvVYNU8nb/qR4vRVyCuCMNjO6fXcMIi5YAt9bhFfoLnQtOdLG8UFA9RLXvt
MCTe/u3DcsXrORWtCrk5hxr0S0seQFQyArv8/MeSJilq1g9gvi6oVN7LcDknI+fvcAREV9YENqr3
F2awKjnGSJ+9g7lGolbAi4sYDNNWkIhHFLqH7F5ko2JpqIUdT5T0iNXJn2oAEk1Wfe5T6dxrpuqJ
ducdEfNLxsGshJ1oRmkf+csBEmDuZdfIG5kiADre6p39f9F+3ERvRxIFKgZJy/PKE+GSRcTjTu5/
e3h0DRC6axtZmZjdSQ3fqWXGXatpAbXyiVhAreTk3q2bFHBbYkIe9N2aEK0ANO7PaBGjQuRxYJB3
PXuEsDGBoFUyggqIjHBIwdyarXjLsT5UD++PolgfWnHOw1NpSjVBiGTTN2qv43QVU7HUk1zC6o3o
d6gh1rU0I0kNW+Rcq2MQ+4Uy7IazgzR+M8KmS6QI5Nz0Mrx638c4I2z4nADW87JArZw67iLh6Hsb
WslLs378IPYlxjTANXsLtnKSd89L9MIqjcQ7MayuIDuvp4zD6ge8tYuW3icXVAwi4N5FaKiTEU5k
AOyXJORZiq3Sq4Xxddb9QFiDSOOAwBf+/DNV8Rb3SWRx9RC2uT/LW24rvTVbQ+w/h66nSbj2H7BR
NNjE0GsA6UepUNbXX1ADiYwpqvDPrtB9RbGY8YG8VwwVO104jcRfHhPWhTZ2TcF4ZjuwiC9j8wi5
sHEWzy0vD6QufuFdkokH3qmX+WmXIVdA4CmE3U6seZuvsh4EXk32ULFNeGqzdyf1F5mfR4bm3JX5
31PeAUMsL9/w+sHdt9hqP3LJbJQkarLJFgIYSKXXu2e9e38A0VuW0NePxeCpMt7KoHKcaBO48SZq
iH0yMzdg9U0r2UEtzR7n9XhTvyNYVBDme0st1hkEdf5nh+F8fAyNd9hraHyILLTqMZV8JKt7dGLf
fFOvUk7gp0vojywFIL7NiCQl0MnpQI4kgns4wlRcqbn7dxPBMMNT0ogaySP7UtEZqlX2m9vmyjTd
CjxxThYhSeNymQkmNjW3mgKCR+OgyTO4r9wtT8KiuNzi1QspvoWJaYsXplmWk2kWv+r2JXXzdIvR
7h/vLJ7AkSPb2n+Z7iZSgbXfPDIw1i8+8T1XLYHZaEkzjJ/XPwmh7O36YJUsTg7TK1mz0ZoKX8nO
PVCSLowXX0BHOq3ZKGsPxdOvKjNXMDEse+DQsK4gPKL68SjeINtg+01sgNeXJMYHt5ynA9F9Wsl6
HY5y8wuYaDg6cJdyS1GMlw72VGYYN7lBhSFx9fFGXyRlCBIjU3HMPOmHcd6NnWpY5ZI5nMHji6hI
UYGWOdrT8LsH61NzQG3/haxB8gsXLnO6fMvEtXMNFJwBI/Gbfn7wi4G3zLIC2gy6Ge6SUXhD+w0K
o7Z9EgnIHpf3f5iB8IIpOq4kzz6QHlEmcNTd81oiZNIpct7wLG3wA+mnp70jyU3QBxafjIA4hVuW
uXdLyzYbm83PZ9t3K7h1p87JGGBepj+4yFmUnCWISlisRdmbA7hanJ6UIXcz5D1CFyXdulIvBomj
RvqRH/2GRGSQyuQLJ9qWOPX1RFuiEGwMDGgz8RJgQ18YdhawSpPxUQ+vl5Grz8hGSXgc4O32zOh8
8+bcDf83RSCYQLUnJUd0V5UJNTydF8Sol3XvoLXH/rR2EKCSWL4vdyxa0TdCrAyW2gIADHrso8VO
WQIEDBXRC3koNcqE/VdCKzs9wr10AD81/LCbaCI7Blx/R+Zmt4fjSkpe+BoKOcC0UTUddY727Zk5
gqXrLcNGQccBx4dL/q1yKGwlDJzLLdc65YbFba5mGNYgn4cfxQYAQDZGwiiEFcvotwU+ncfdAZ3g
udv3nIo3eJbAU9PozOlgNUiihO45R1VOBgP6qBWVWbJt8+pKHG9bR92RtI17P+ssmqUbKSPBrOof
4MOVr0WOQh6NUyGwD7X3NRPUjqENMbWKKWzmyeYPQ7dRuZdm+TmOpwV1QGenirHXlhoSxJaVu4/a
Dt0Hktsf96hmzj+QuqWF0F6n1Om3By+9w8MJjbCoR61LGm/St2EsFrZMHhm38d2U6DRFe9I2Ajhe
te39GbddE2Pf9CoH9oYW2g0mkc4vhpS/Q6Zd/pwKgesVVJ6dghVIKgcpPV3qR2Jqicl1cabxkq6D
r3+cIZCybvXNhgZiXY620giSbsBxgdzsIYqnKM0wdDwrXtp1v8sxdPFFk7aT3tUnOyOrymZtnmNZ
le6INEMNrGbbT9aG32bK2O4m9a1TZWB/Fsk4bgLHqDfeGzGczvpByFs858AQENXo4ymJ8s9zWy/B
CKMEKNMu8pnFMsOdeC81I1RU38llkVltUgUO2ZDmvKnlSKTn89XyKWGn3zKbaTuFQyycVC68/ZPI
FGN7L1eEovfaJCYRH1DjqPdxlLappevtu4Q2kAZmm29Wm+idQxIrvll0Zn4hWDCAieesV0LeOeS9
My09FTv7UalhK4p8uucltUiMfOG0GSvaDjpdDCdbIijZSk9zr4edf3oxxel8n5XttpkvWRZ0Qh/Z
ZHx2mJv/t0ghzCnrsu1TDIKXT0v7Z9yU1i5RB/yRnwa2xO7EL+47eeHzYvafB4Awj1hnyhbgfG7T
QEZ+P5G8ON+6VE1aIk8DtvpoXPJsPRsXupK3dfN/CffDeUgoB9ONNIek0cX2c7EJOiRlyKeog3Ou
UlNni4uyO8RZhjAHZy7d5p5vBuhBW1ieRwlcR7vnR1hfbf0iPPSlOqq3k48EZ2V+eG+us6rbIddq
vLKMoCVJ3jP/9o8iq1220Wf0yC2CJYvDdUpZIY2RAyMcefLLkPzICxTRTh8RnxY1RFDcQfr9WAnE
agYzhnAgCDogST34cZFNQNQ++xg70zH04I23yTJrBrP/aSMpq5g582bjpGoa/IHwWg9qBc48s53x
O1NQTnIvtld8n/nn/3+t2szi2XfbmTYwReLrpcNnGUYC/v6vcS+7CTsJ2MDJr5o2Y42kPgFo8ydj
cLfHLR1RT8UTIHFvj2X0VJHlJJM4RQ7bBsZ/ucaJPuJBJE6M4HGUO9vdon9LCPQsShOUbrBLlK4k
tmMFZApX4LFhNfaWx5QkevG2xH9C4Ctn2h/YGO35/6Bmb/SJ5Y5+OPFB6/TrsJYy3401MRVtzp8p
kmu8qVOGh8q99Xeygn0ha8BCGINFWfufvPKPmwO9m04upvy3WpUpVXD12nA1Fsq2wwIzaHaQQOwF
bNHWifWRE5cEp8Zo5fack1ggCJuPJNdKC3YUhveEDPqYJMIh+Dv19InVCJGt+MI0+SUvGx0wX5h3
2U+0OplWQO9UrPpd3NINDqYEOJIi7IzvpkI1wuRiYZKXJg9ZyoXUUyfIYNd4KTRhoRGXhuAU8/yv
bwLPrbr7A8kwwhSt4lA3ddwrw6OmJGGakaDutvrxey6aZ20hJqPKGSXsO7ky9p0T9jrXYtg89QPK
iyo+9mRP1UU4mpPQ9fUcFgf0RNSV5pEXDJCFmvI2iPA8kdUuD45L4bDR+rcBfYs66gYDzgGohMXc
9j6BFqpncli9fDCOddRh3vvBfJlCyRT1RUwHI2lNdkjK/B8Gzv1Pdp2hZOhRTArusxrKQ4jxzHjC
rzcAqS69jU8X+ETusmbP6+UDgAlOq32I632xDVVVPy2MetbEwdntCfSEDxQUt+24S1lmZEBSyu0U
i6ybZJ/6WsfC9/5xAxA468Jv2crLxmzUOqJzEC5TDSgM0iYzmG+K8Ect5Br4RJdBwbo+ccBuhnKl
rN/UK0Waa4svhfgANGvWYjKa9OF9TUh3HLZ7N7+ssLQpChw1Qj3DNbXq1JUjluJz/iam21pZrk/9
LF/8yxxeazXWsVkzrP/bwH0DirYVbYRRq/tRoEr4ys0qOOPb1Bv91EAFZGxlbpamqWfjBlnpcyL8
EoF6yI9rwB5jwHbsCRQ5W8lMfv7sKZTqseeu6jKteFV7Ei2BbqHr/mYE3bh9biX4fCOL3N1bGJoD
qF/ehb2dQsjdqOPjOZk/FM/fq8THxbm4WKq0BY8+L5F44GPl1wrsDgbUcLI2Osmfnj6iYJo446/d
eEKvyW3DbkvPXTDCHaEEuv8ZzdiwOH7xw5YqYOZJQHVm7t0X5GQmXgXB2/wwtzuM9aP8hs7PELTj
vmt1sMQumme2F8ea6dcWlUaKSjMOQNDzWyUOJwEMHrK0Uyp4x0sGIZYNOB7Q7d2U/4RQdZBH3PX+
w+v3AoVPqORc7WtaWBZynMSBFYpLWlpsUNK13kzeklydMqe/KEU21aUzAv9hp0SQ1r3BAfY2+WS8
MynW0OzZPOg7YDximTaa3ZBVTOHyEg8/Movj1x3ouDz8bOAPoP15wVQpU8Csa1ESYXGc00y+Zttk
tGpt1UE0ZNOI+vvlVSmfwHcyX0YQmDN6TEsVS89zgCWO57byELjK50gIc41ZkV5G76rvkbZG6Qz8
OIJhQlul01nkQiiSg8NuPMFJj5jmfQU1fIyiQOeOExaQx81WuwM5d5Bc7uJ902ReiTnrih8BZY5D
t2x4EbXfOnv+XLXrzBeAdpVMxE5L6WBNDjZMaGjKrHgxM910eMJ73FUuT46gnEoxT4Z5Wg4nezRR
0Ftf1DVCYwesQa2Q+kt3tREmQ+gjjHDYUWJQMeZEcc5+rNEcIrMrnZxuwoTqzvk3dExgcWwOerqh
vjtbK1xg9b4pAvFTy50lDXeEZ4vuA+d2ZkpOKn27KKEek2cTm5hvTqKRMhA7nOnRp4nABE4WRef+
2NwHvC++B0HjM9gmax4ibENaGuPWchm8BJVNrZn12AJ8KCZ8qA1kHS3K9KpvGKZIRbwfXf46NZxo
A+AAuKHq7pRBJe8WXU4cnxsEalzCadiBd36JWJaZOO0+JPeqU5YzvufavnHjZ/+zbuk6D0To+tOm
wx1BRp6E2R02v5Kf8T66u2HT2axWg6+0TO3Su22rDhbwx165OTgE8vp0iGG/sBONNU/w4/TwE1In
oZImdjNa94j+qljEfeBeAzSgamTkGu/veeuCk1FxcxoN1Gwrp9/wYb+sIrdjgx1mjfOgl1MKoo/5
ZF/djdkMntXu40hdRmWo47QdArOgtkP+z07Jm0ZOfRmp7akSKKr9JzMllGSQZ4Wzuinkh17JnVb4
bbfobtcFvjM/FNhMPSFfgbFzXgBEmsTjn+uhZThi5UCDk8cKonF7yc9Vmqk/VESqyZloieovC4Wp
InnktOje8K9c0xGS3HPoLMHHMPiaGPSkGpH616EgUZQnjxvIKk9jyRRYmKLuB+yB1Xnn9kQuyEUK
trv6KWdhyRKoalRw+NQ2NK4OZURsCrAGGK1A85d65Hr/DvJHLgMWh3aAqshHx6oaNNJxm0FztISO
E7io3IPSIzy9wJG81jXB5/RlpgMHce6DsmQKLFEbdUS8CI73gmkGM7UhT57cFpGvKx5qcVm9dKl4
scQo7sjdFF0D6fa137nxegIAzFP8IuvlSrO+uRukIk0Ew8zefRuFk+5OFdHwqyg5Iyx/50SwlNme
1phtCDln7CTrzLo6wzXmmMBmGGHyambETT+Io+WTo5mJX/MWZ78mHw9Hot0clioH6tjvWy6Vuww4
afjWE3K1SNWqwFCncqnVDToo5bLKZBsp/kYroUne/HgmJ0PsX+p0B06J+DCg3fYXQwC/ZY4u41L5
27wzBr8aAyeZkoyMg3I64he8C4ZZx9uawpuDzf1+wadNUna4JXuJfVVV5qB1VnDW/qd2ErCv4WXy
oWilEzPpvPxqYSmuhkZolQ1B05lNP3JPD9uu0LrOfES+4uTO0v6eDaBD9GVjkry4+1acetUxs0V9
kdDrHO5L3B1b53qUF2ylpqCsY3tJOdGDOaVzSt9Dz5PTiZcSBN3HMGLF7cx1vMrn27uOhYqa+486
LHE+7Abs6lU9hagmjMrmVQp6hFp5XRbAOXF48Xh2F2z1M9bR6e5UWr6iMxAVFUBySk3MPqCzNKeW
P1Zdz86a/w1Dio5csvnbkoXKS+R2vZZn+qv//83NOrPF5xA3mN9cF5IFjWgAjbvOXHIhOqZPblmK
wsYk54FFcD1/Z75bz67j5ZFJglyXwc61RAw1m0U/wk40VCJz3idFlw6STT37D0Lq9RdmohajmsFd
Ok7I/OrdqiuR0MML03xT/goL7Z6nS4z2uHJyEqhWr7lHNNKwap/3woTkwJgU4zXeMZcW5jsaNHQt
OgHvVh95N9z00wpeCCnx/Hj+WRAY/r7oafdELtpSC93vWatp8Sb0LTZXI9tiv5wew9qJHNM9k/QN
6osLYlPAxc6I22zzM1hBdKLW9pPnmy3hGsLn2ek+MsqxSNuTgOXRow7i8o+oT4kDd+5pSW9QzGP0
5JGfJzXzun3TZffdL876D0SksmAJ/qqWXQERXCIe2r9udaTpic+ugLK9wIeCyK73ZOIXb05Iz+DQ
00r+6FRS0EFN+7YSfS5ArTIazNuFlc7+tGCfTEIoNAYTgebLkCsx0a285vBXXBLXMEo1w84eK1zT
1JDXUlePb386iIOCe701OiBz9lTJwlmn3MWN4r08RKF0Ps/1nvwnHpsIBSrGdQYvfSpyjrt6+Qt0
hRAIlpbxVASZUdOzDj+525vpIig1jTNh2imJiUs6YkF2dCVLUoiXY5IHfURnDSLJgaHyGG0QCUEi
ecEsyeiPcZEg+jbgob01ydQljdbnm757BDooPQ1RlJ9g4YTdnRALEkewlvz2zjinEzttA4i2BZ8i
uEqgxCHlM9uYn6ebJ9hZyWf0ljqAJt+zPnmvouMvyg2IocA9DpJ4MziuI8ewKsBVW6Q/EfAha/5w
G1iuzhuw7XdfNYcx3kNTethrhD+aZjy1q7fF/7YViyp5oyz3tfRSmf78Vg1OAFdOT2vF021SMApi
NcS38Px1tClszK43V5OyR0qiKR1+l2XcVlgw6jnTla+Sje2iC/L5yVIcnZpBbgPSTusd1sS/QJZv
4Dy68L83927w97MH9KwMFEZvJgmbDl8Wr+VKcKHgRowb84vv1lyJbSDAKVXRr93Lh457O5EkUjZF
IfqqXuAEEIl4LxgANnmkFPH92D+Ialb/CEqNxtgiNFA+4QZQlCYZXksG2qgENZzU3IzYQyTRn7M7
P+LGJTKaGJhw2sdPNa8aSY5aKV6/Fg4EQdjGisJHGomJQA0xEYyd2SEk7Eu6jP3QEZU1JPmvb10K
NIsn4NEK7Atp04F8HECmpboYNCyUVRbe5MJhXUlmWeBPFze0oSLfUtmPWHNZVr8AEA6MABheFqqp
TJyagITrAgGteryRgXMdK3mQK2Kl02mk8E6TiEu9h1Cig8+3nJDLjnCCZfPka9fQ624HVseosyNe
Zqcf4Ey4o6/p2gSxQt1niyqO2qTmvRjigVeMF0CcKVKxPXFUs+h/od299qUBFLG1/yhFjr66CrEx
7ejq3igZ2bCdomRG8P0Tr7IC0cKVaisJ+jgHFNjImRUJVu/t0k0Ctz5fIwtj501ckjho7Q5VfHgx
7EHCUIDmHCRVnKJxcsRVNzLv3sXJhswlQXr4DRqQmxuCHLX1Sj+v+Ytitf1PVe60bDUVw/nvWnid
kwr1vVwhyoFbGCl/THeBM//l2ZBRxaRPCNDbOktCkuGBZoadn9TAthiJILSLLLX0OuHu2m56gBx1
rdJjxeGfJfXVGjlb3hEfnDtILnq0wo40Ou9M3DrIKr9MSeaDxI9Ow1LFqSSWvsHhcW6jeRdC+kzs
3Z1eTpHP8bk2hnxVPTXkcGI/1dseYSvHKXQR/qmMD7ppnXUrIPRClr2G30k3vl18t/DHechr1ewu
mCUhVe/hR+Jfa7BAcxeCxgh1E/UMWNzEFWyDLhesQrvEvzjtDoJIPHw8V/6denJOtD3AYihSC1B3
blt7qEZtgWYMbJYFKjExU/Zq730SWMFMrV1Fgy+c5PWTuvhyhEtOQR6pTscyvAttf3FXZmpkXQY3
kdlKpLpjAqRQ8Iu9EV+GuV+N7Zk3th9CQgjcilMFrSAdqK8wOhLu0VBw/cTJQohRt+/cNw6sJ7pD
wtXar5bHDQTOrN8z/CDSl8gbOYjFQa+VykeMJvhc/BfrsLg3qnNFSQ9xuo7IPUdzjNvnq1JhA9y0
xANU+2CE1pzCPpp6O0gsuJUpx+DKwIF+WeREhAgCNGtknLzKlrTUU6GT58yeDKgBdXfWubhrrz7L
JFeCHo3f3p0cCfOfbSfIIYjfS74aAQpT0DJ+Yt2jpak5cGlTz+6IgjikaUU4Kfb8++qmP20NX7At
3Bo8IgoxPJuCzzPBNmSZk1QiXszCw5Up1KsLCP5eE446GgDe+y45ldoSJ9K2+8+M+bUwVkz9vyuG
3YSqYolOEbIpLQrHN5f3rrPV3AdHUmomd4FziC7b2b10CSKVzCc5RHEw+1MYxZ8SyaBg0fgWp3qb
EnBLKXx5oLppOJktZbcXM3mjFh6oIr6uPFJIR+/0qhIy+LB2G4TGlwyHKpGUIL7gpd4BvrsWRWQo
dDuIaFz6V5WTXTm03OrcjXJdgoKmdwqcyUFV3bRorNDrJ/SUDH1o6bNUjOFo7Tl0kKKAxXUZCNFA
g6kw8MZrY5gvFzlgMzX3B6t6jpYaZJKxN9MVA2zmgEraF0KID5MHiFGY6nilg3tPlwpbPGGPG0sy
3grwk6VakVin/BcIbSrRThs/4Q97b66j6w5nSskEji7WZ1V8kXbjNLnchizNkIMvjGUvf+41CkUy
COqiHAMunj7/eCYFqgri9MOvIOXh198fQodwsvYcbVVCheUSxVu/Mjsk6rWDbXDdCUsALOVNiHYI
YTkI/+arcCZPSpx83DKVs2NmIQ9p6itORIH865OP7b2h5VQ8u+UcrGom5FCSJW4qTZ5o8uuxqGPH
3LJ8h65ExcE8ARHVMoL/Uxb4IKcdjtfR1NlQsfFkacVbZyPZ6B1grvKnqLF3JQmmEo+uHcNOJHfL
N1nfE4yYrgwc5nFhHY1yEKb6ZCksCX64F+Q1islO41GrLGKGW9ybddoAqQ5FGeNiMHWnAfGMiote
ujtpBp3UPMSIrT3Zj7o9OvNv4N5ugQMjJtk88PCFpi9nBn+6/mU15FzzAVBi7qu9TjNHL1Nvl/d8
fnHifpOwE43236AK3j9U6oDJwCOMiuXSFd93wy+9RVikcsmaBoLM5DLumf5JVQoB2AVcB+Oi4bH5
xN6Fz1GZ6cw0ADXst8Lpu4F7SXPJ8u52mhHnkojA6O2p2oqV9yZtL7y7l3cOaCo1Hqdsmqa2/SCP
C+EEvdNKn1MkivfzRpMJxo1ZhUraMpEZgoW+ZxyV9B4FKOm02xhkxBU/frvPliTYcbHjEck8fqGX
tZ+7HIPUyoYwZYpPMX5aoovOh8ULGtpJpIrW+6FHHPMbtmvTTM3JmgUT+PUOkoKip8ETEeHmvZ7G
kfLAJInjVGIm/b7qVIbwM4a9L4b0pPnK8suz9fHJkwFa/bZ03pVK3k5JYGJWI3zuSvTbaKmofhOz
9V5JGzToE46kYiCCwYLQcAtMEMN9LwA2/ZJNBj/B/gdrU974YHP6w7BecB1VolficDM8KKCTy7Cp
/qBy5Cd4rm7L2C63c8/ERrQLX7c2pFCZ9ZTnNPfHrkC1M7p+DzRmJZPpWjAqXF5EAlPfsRCxSPjT
vBDiFMPW52rpNwPVm6DtVNW5jzkK8hU6DwKINbEBEF16bwdh/u0409aApLpt/P7OLWvBuxE//sg0
WL5parGnhSMRTdddKEheUkSwDhaawrsU4npq56COJ0jawU3dY3sVDf4Y/wut69m3LXyDvKd8Vi0k
1PmVVjurh3xWuBRUN2wSE38EXCV2IHeqK4LccQnayEiv/Klh4dMMq//3q6aYB4BtM9vEZaZW09c/
4n4PFQ+yqkCOzVfw8eGQYcej/1EwbGpbvvLq+4Ed1VEESIR4BsOO7hASc3IrQpEvVi+u7eUnygf3
4hm3OK6ZDX+SFY8OJm0qplvRxXwSyKJkUFfWGiSOQy16ZiOKnuGrWZFX4AGijkTEzCa6/NGjp1kW
E1/2GukCR46gXQ6Xcy1GJIJcCTG0YUbmLIN5/civVi49pLS+Tp2Vsd7Bx0Qmm19qCTl1NlURoPHW
Nc3IcSvUDt3zKM8FbLM5ZMl/OTHpRIaFXTPXeBOgKN4rcOdhYSRTYD0vVtfCQzzHyUl19c994/4p
LJVvlLX440xChpx2mgRy4NN0bdf0fRfUNGRgoptZtshJ8tId4zwDdM2R3QolnOXwA6Yb02Z/6KT5
ER612dEGyBlR8DjfRglVLdcz++DKbdIc3c3DmktypMkrrNFt06y5Av9Re/QO/ul+6Rh8xaHJT3Me
zj5pppgdLYUmeCTSSp6VO5U0/xw8DH+BOHT0nAMfGQ+9rg1/zLvE/SFzLFPsLphYtaynOnkW+Ktq
EByypEbMYdytFbhILv243n1KeOzL6bnFgn1J/rJPCOXWR4zQPHh4PZPRxWPF8jtwCWOeQldtOlfE
NJyDkaj3xRuALgfAqDrf9tsBBftYLX2uMcYt3Gt+ysOjp4tIE/rbrMW7oORg3ITvw0hxflkGSPU4
KEC3p1d5Npv4MYxQBFT9Xrp/Gx9ZW5DRFmvewg22O2eOdTDl0476MPm1E99hm/91LhELIlYqCbEx
o0IQ/fygfWOlT9uIGAbnPYcsZZvMtfb9OHJ5kn4mJgB9JpT8vEXc2XrcizeD3FFPdYQtaYwBkB5/
fzjSa/1+wkjCkYWquXl6wErBU8jInapFIWJgxUvZUwZLuOmaUYkHX6tMde2WwZqtOulzLumqrMYQ
0cA/3lNQASqEIwshf8+ojxLj6MKyTOe/3faO+uLr1lsb1Nm/8uBxtkCjHfhqU8YBiEn9uYch2jET
iynYaOXpcDAi1JL108ks8lzGmt8t0Pvxkh6dq4ibzT071pGUEQ4hgusY/dheRnPNVaKWFKemOkNW
S6xCpdBKWJvHVv0onVquewmaHij6qk6nTHaV4gITTUVJbZxjeDxUEvWeVyOpk4VsSbsxyvFDdNqu
mWfcd90A29cxrLxk8GTGxDOydcXFMM4tKCnuQFogqCRnBKxKXifHTzPccoASiWPoDvjwE89E89j+
tuRzn2ZktD7pd54MQ8TVjjcqgS0cic0VB+IrQvcIWqBbLn/Wei/P+uG9xppMRpMILmrU0WLIDtNT
qsdCF2HI8PwaBEMctwOwIiu1MODI5EyRJg/qK8Qgz9BjuVhwdHZoa79iZswgBbg0BKLyzet740m1
boBiQCHy9+Gj+ku06EoBYwX+UfG7zyoqnVqOGBqoBHiI/9EbaaswkCoPqlijBfHYzEuN8MMTBm/b
3iTEzbQVQXMEZ2I4WYE5TMxKV03+J3NeY434S3HPyE5S1TxY/I3/POKaTrfFwWfAJNPFP1J4dClM
ffavj8XJu7d1eAVx+tSNpsnXBazPIiGxx7QUziMGjsqssrvxCAVSOn2DMGXhILRHojUd9L2hV2TB
zm+STCPEP3f98cGv9UryYcNczQp64J1z2NJkhHaodVFz22WqODiwFYD4n6CPP2E5BIPEYNVNNALc
B6aGCtdQbRuKNc2zpuTzhdAjqbZ6C+4HTIw/JA5Was5tzbOKnGBX4LFJYbHPnG4hwMrko49utAap
IkKC5tel4ZmisexStaVLh34rCDmA1B0L6c8VMvLu37OL8Ltd5/5jHiFRa8tu+v3YAl9ip1dhNedI
N6u3SbsctMhSZhg0DYNLOle5A+6KGqUfP+m82NhEBVGqC6aQosvtOblqMpnNvCuhAHZQqVMl0Sh8
whQyOmZZXxWIaLv2wuWrB+NTyO+kASfEeFQq37YFbWGihDEB/Bq7sUp7iIzCYkjHGo6ykqzTBBvC
YtYcQar3y//IiHWMatDVsoqpiWDJ+iRa0OpYtjEoSF/989ffV78a8mkjfeah9L4csG1yTSieC05W
pm01fxxMTHXXiF7gDfBF4dD5+RNSQmd5P6XbLqIGwF+UnhdB9FUtF+3hcQEInfDEA7qIQ2bDzKOi
bmRLxMYuqEsYe91e0hA5H9hB/mCX6BTMp2FZzx7ozTkdGmyb37DCemFbVmMb89IE9OiHceQ9Cv20
tiAXQ47vDaHd/GzvIidche/+6vjOBMy8VRYtL0duwGPlSBAIynaLttaewSolTx72YPo6UPIM1jh6
s5BETOqR/VUkzPFtlkuth3kDSvIUBQZRqm5W/VP2KRTEL9FGXLZhHxx/rl4YPPVDiEzqJLn48/bt
/f9mlbg1WePf49awOaaHGhzgILEk5x82IMXGODAcuXHOJf3V9LYa7cEOvRYztPDYzs92XmV2h2lR
taVtrUI5RNtb5BsxXttI76FkGHxX0fdCRi+SfDVMvlO1svnHux6LlryXzW5I9PvdPLJmWDG/hYWn
u6RYDn52M3U8TN1GrR6c7cBaDlpZgxRnYj3vgQRZd9cq7Hizme+0LILzuCX11kxo7pQQmfuUxYR5
M1w9bXSP4GaElEo+C08082PuhPb00ONrF9NiYbUZE1t2g+rJ0WZNXujIX35KbBckkVhXlOf1ug+1
4mq4wVbz93BrVnIvpMvW6CcGqSASyjwUXcLoZkvu93lHZr3oUthyiQ6rtRe+KVrbmZuiGCoP+wKy
CjJpUKACjEFiB6CEPkcQSFRa5khajck/oqpKtFtMVN2byk1YorrC85Jx2jx57VnuY3D19DUE/J+C
g5qyoVBzbQBaQltOlAQ0T6osS9ocGF9to8QglvTLWDwaACUz+sI80L2nzIsbtlUxuEzpddTOoS1E
ETT+mio/e4fEbOTbfq+HbDZZSRdNTTwdDoWD3P7HscaDLIWVamSgcAsLCMp7WouWUJ3cZdHsADq8
vd00rQSD3BCLiYVjUbElXv8zfWK8WpMPpnOLesxiJxezuQuQ4ATzu6gojQl1AfIaTX77cd73Eaj4
bnnHyZz55ZRFYwXu+MozF2zIhrZvuu9h2nYAxJz04cLGaD+LgKm48N+Pamq13hZcHuoMFYZKvcZV
mnO9lIak6FrFPTNfFH/Sbn/QItinTOzd3q6GmJKWBkJBEqt7DFr7OO44nSgzNXl+z2y8p/eRWnkI
0qr4lQAAwkQZ8AqI2gLMs8XUIoc9E17mURRLXa/pzhlTZJIzI3qirh4tPeMp+7sXVVyMo3mDiEK2
EXWduxPkAiObLMsfhYk10Ciqjwyg8W5ERhB3hqYJNj6avyYOtjmJ7E6hwAnl3fUMZHvrlsapsZc6
ch+CirxzSoPUhS//ZButfCI2VQ9sBGXaQXCNyTg2JnGnsx/xLjvaDrxGX5Nraho0WVnnHEFF5+Fu
x1JwWktGCIATAJwFLXSuCMDG5xKn7WIOBVqYASwQwyMZ9p4GMEMo5kKCI1FOLDUyTpYV9ZrO4YZj
um8+1Dl5Z+uVQ5bh6lcNOeOvSTdwoI7XCCh22RTD5qUJp4WE/JFqOR+ta24NHoZpS3FGYAPHN2Rq
Mu4drtm0d/3VKcmtVwB7B9hMLBeHKeyjmHcZfzEPA034EWSQYyYc859h6drK6w71V4LnbWRCLSmR
MpU8htHlChUaPNjKYWSU9mjaUbYg4OU1c+sF7zQidTWp6jYRqmT+qh+3vqPkS2XxA5j7qCBO61vh
sTgqKcKLgcuOLD8XzVI4J2RC9YiFFazbj0htgdnJ1vqldUVQx6nJ5FRqwqz8s/mFYw0eNakJ0t99
eCS39ag1efK62qvCmJEzBvm51WEW93Ay499d+tMjDjU7O7YA65eCNKCQuULhZCeymkh+Wbm1HYwp
yFflcHEqZB2YyNZmscFNBt2qAHyPgSRvsvxVY6Z22+JHiS21ytc2gJ/8ZrhSd8tOimKuboPj8O/m
KFSvonKXgQorZOPlF80x2vygL9T9uzMxcNQnBbS8fVVbFanPJPVHcMsKV/KrzaAVIuBcV3TwBbBp
Zkgflnj7G0nKfrWau7ZTYdc2TzwaYanZwimcMcvStarYQEhhWJCOouTBtv3k8YfRgHrTvzaZfFZ4
51ZZD/+SzdKvztiJNaK1NG5Xk42N9fC3LQHHEnhU9RIHGgWgt2BLeUcOEnVEA/x0AT71RC/IBa+B
GICSMP4abBy8RDU32K/Pe6kkDpMhwn8Qu5CpUkearMiKyoZ3DMp1Yiy4VfDEXYiC4UepBGeEo8ha
ybC3STp2LmluP+tlFJW0PoiaJntMo08igRF94mTXAHnzmICSxHz1GvnKclEnpfzug/nzb1gnyCA+
t7HXFs/Rc8O2kXcErn/GeFW9OokERtO2A0NvIcpXBImDxIHo+NZVSLb+kJhc3nHEe9l/oh9FhFEj
Bfdbr0kPmSOMxcnCl7mphunoJRk1Zr60kpBL0UZqseWJwcEZs03sjeXafPWT9wZQDISUOJDJn3mh
9m0YNyvLMgv4DCQIWBcULR9OU/qCM5GqL/u3kUOeQk1m420mEx5V82Iygn1yPwoYYWj7RFBmeXV7
W3XGywg2xXjMbejCYOf+PyKQOC2doSy9t5yG9LGuaVABR+zk4sKCHcYLGV1rwbEIUGS1fcGo7gbf
7QfzoXWnvxpilQoS8casbRxvc/JkWYzWGRxq+ESuNhB360wEzLSW1/0GocF15BAuPK2hH1ABcsqK
TSFljThHv5oD5UVTuJUhoch6W6HDz5FDilru3P6G6o+hWFyaZejg5DVlkGp7tbvLV1G+WZR4ZEo7
aYIgqkDZOkYkHWVWhEilFwFxf9lkj3qKB3AQXHVbS7A8j0NHYxwJ1DqahN1chZEHWKXH8BXKrOXr
HEYzwIGoF1cfa/CzDIwPc947RUijkcy2QJsfEkchpWGhmgQEFdrYpXt3ecraTgHKPSF9DRTxnyKf
M08yOVUZGBo266BcozUTnbugCVUujdjK02GLTO6SXRrCeJwTaxJ63VEs/bGu+MIxd5h64UhSgMcN
btHOETj/J38RqQU8QTr6/ML/j/xH+2Kq2Yl6lV/SMR/nO7rLvQhBS/+ZNNwzqrbNgYrzy9Q/slpP
5QoFtgnsoaWGOI83l53O5GFbAyAg2NWQkNphS8lk3hYO40ZGOF9zxyCT0nLp4YwcgewiEqpv4Iug
PzoTnsgT3QkTgjGew1UsPN0K9xyvxOgyVJr674urRDNPlI2vu+Y/5IqXmPEGd/jQfHCVfk9EMnNp
2McyBxM6VZ6YDMi9tn4r3duBkJ0TEXXnE+1I6u9LSBpgxxCGH3gKbNutS0Ai7VMR26iTEa+ycOSW
8dg0gNygKSK24I2PaLIZelMRSd2FaPQoTxebUW8ZFz4PTj4CnVdFBUi6K6dSx6nw2vDTJ3HkygdE
5Ayn1DoAhhbl9hZOJPQa0wN/ufoSNn34r5RHY/z1m+5+w4LJXKrhq3A83ct13SvjlAcDqrEl207Z
6EVLrmSStOyBdmXmImvmeNKUHUbNSWTcgIadWECuI5RrL/TPGKbmb3o0C5cznzuluGrq94wZgBl6
CYm6GqJufaSAbCJuUO1fCBkztI0/hK0BxONM1Ariq/oXryiocI0yjWL647oCotIjJ67EGr/0vVb/
YQFNAYxpq5WckxTiqLZ+z+Cavsq5Yoop88AovZ3GssXO+GtoBmouA3Eqpsna0CKXLaSg8HMSNEXm
8wTjBEpwaP/PpuKaTZOxyc8ew7wco3yb4dwhhFzVYN286ElCRfj5KylDk9rmCIoGn/bCIOW02g3W
3/ruI4s52PuhXXwkrEJWVCVueGj+BqYbu2FK/k9mwB1Ft70OZQ7RyeklOm1lwNRAhw9mqnrMmwB7
rrW6DwG0kbXhM9RO/1ibvWd08TvE4GvFJ8+TfxClUZMkuLG3y55QatbyAThbHLdYft/LTSUjR5PO
4r7Y4y9fPFpVveRPIK7joGUO31zEenHwCNRMtaQ5OW7L9Gn08rzKosI4vfFhS08QDrYFGcdSsc5J
ffNhCrMrjw9PUYgOO3eEVYBV7YSUo/TzSfH610t7VaoblryyYC5PfKVCnxJsncJlmNeQpFyo7rxF
CMYx02dx9GuVYQr0fLvaaF+NhH4sOAW3dCwSRlq8sgoLWHCqxODDA6pkNV+ZMEnzQGhrA8yPrxce
+rK60PVI+/lkHL4d9NWMwxu+gdsmNfjU+Cni8Ay6M3TIRkcES3y/cIMmUTQcHpE84vFz/VBTmAwA
cHjtSHTnbWzcDWatRGvUFSrUZh5PL2R3X3p+HJXQKpGRl7b+rOTZgwwZT2kueFxlsHRNsFzmJKtR
9cLu+kFX3gsiJGH3AKXe6QYSRUbEaFJG3fpUxaYNrPNd/fXRSQVux9EgzD9rOZFhz5Lhv7TCevhS
sJNL3ts5sC3CYp5HqBzYGKqOyCmisTyiWriYh8RHPqJoTQnGj3BP4ZJxe/w7OjmdE5WMYZ7KYlcJ
40yOpLOVdLGPPjLUZUYNvikCV5bcBHVvaLAgE9BZwOFFd1d6/HO5OjqYnFQAqagyUZU7IY5jC3qx
LqVr0zzXYTHepklqShMNedxgD8nHE2VhuD53jppO0pHIp3w0a3673OeukCyzb4LrYWgPHzezlanQ
JWyVCIkgGL94hXE/blWoQ/W4UVspqFzKMAqAK24PACfzfzzy4tZMFgtqfTgVnaRD893J5S+V3bMa
Gx2f9GaC0jgjOnb2xsESdIZ31IS6jyZu1SjYH/cYXeC8KzNkL+x8ZJ6IMIh6862KVSWna3yRIa01
CFRM082FpANG2Tpp2XMPtH6WuqJOlqwoO1QMZ9yC6anuuakUL25sH1OCEU9gmLW3y5pet06ox97O
BtlGiJKI45xjIkGSY7u+BrFYmwMmg5PkWZCu0BVMTe8mFFt50eF+D0CzNLuGzRtngz8g0GySc4Za
w0dTy974MY/eRY1AGYa4eodapq8Sd/1cTwfDaTqE1GcgdsVmIzU64H6WYevJIe8vrFW902uv0B0K
R1jar2++XkXDFe7xESesulBNat2NBIAnBrg3dr4CQjEAGTX+PKq+Z5oy0zpQ7J488tJy5BqkdhY4
wAp5DwfPWkkeC09TvqIEwST3qBC7gxc75iXNdfllwRkIpYCd6WRiAlHS6clg8Sbr3jVWtyWTNDEr
28bbshJzmQNZjAjpbFopLGnsEbGw5gZqjnR9S9ayUI3azx4vbEhCqiT/Y64ImwSlqC65wTP5ZDCw
drHmngfsz1rmwku1E3536ITINQY7Lkppz4h/FaG17LqOi4dv/gZG8phxKmDlixCMYg9Qxsx8iTwp
vcIsXYwt97VAnc8dD/A9O7eRJRreCXecTRp4lgPNVg3x4W0aQH0CMIa7paPwOiwjJUBSkbtNMyJx
zXcClytdiKoSr5Hou8flslW9rCEQt0cmX6dpS94zsZ0qkePwzDAa+8y9MCOU3/shZOL7dYa4bRML
PsEpz29fg15zVIl89qePBEsz2HUKTP0dT4y2v5Q0AIGs3VefUTZiU+YNHRXPsfugH8l8w3qFQTQg
TK7iiZkuXcZqK6GiAwu1iMiMhoV+Nj592EMZh3UPBQWdJIx9ktAM9Yggl+YM/EG4iSjRAgALy8MY
JBeLZEAzKLHXYF9aV9LKcqAD5ML62xLPnYd+411vZBG1QsnqoorL7nUZE27SbMzD0ZCS8uEcNsPg
hcrKtKs4v2GQZujNpHlMtLvKjgFpUC+2d6VMc4UxdmqoLlOTMESEtSFJbltZ9Pm+xbgrBG5jv7Sd
v4HnFtOS8K6+9EsiMQ0+U2b7TdnLn/AkgPVtQZTstSXxFNtOWNFcfYFCSkjcPyUklX6czmHd7JPv
Y6E1xD9fQOPmgPMxlnvBJf92iaynu8T5vncM8Jx/8crw7VqwoTsCE/FX2GhmVPIulgxBIcbsqEL/
7gI81LpuU53lUsj6HlXb0FFDwx40sEQg2m+7ozhAizwxh/OW3WcGwkxtpYErrvxA0+EWtFfCp4Yp
8WbYAhLIpKPVfwHNopebM1OC7ct2EIVojkBx6ZcnGLkL1xPJKO5cU0FkCChtiKNtcT9C+adF1Ybz
V7hI7dbWcjSHNAFY0Qnf308nNuag+z4q/S0PBNwctOAUWn2ljIcEbqheghfWKwrq2EQCea80O891
XjSxzc1mfBi5oubTyg6RZfQ9RkMT8EEMuA1xoHx4FA3Xa8Ms4ybxBIMNq1EwQiOwyY8wqE1Srvvk
/ZNpEPgXvZOkl51GnbnBEaEuprW8Iq6acAj4u1glnYXFL7DyvAgziyGs8YNEx/FSSn6MJtqjt2Sg
BW261Sc36fOMD0Ub8yp8nCY6F1Y8+VFSpmDO59qhBbqw5qWRwx02OfQpf2HVPKnqVinzSPj5vcKn
pJ8twdnMGFMDZv77l0OX/ICsJz02YTtDEhvt8hl9lnV8cGFfotzrNl/ffsYgSnBFEVDdCt1sqhKQ
LaPbU5u72rZ5Xq7EMkJw2ZqD6o9YlEGe+8mOi7YppJ8mG1NdsEJmDnVDKtuBP9tCOwUdORm/vSIK
9Pu3notI9iNc8uLI3AI4t6mmKWcTOogLTdU5dbDdWYVtOyoDR8ak2nvoXrDQL63YnDkhbiF/So0j
/dTBulVp6rIDTpCJ76oINsrKe86dLSJ5rCSn7VHGqlawFlpO8BwevdOoiviw7gXD7Jkk9T83WBdk
Q057ejlItX7RXtd8axBG0itGAyqOGmLq33GNotuLh+KviRFO5zYZw+CJmB0z2GZY0ehM27m80NMP
vVQKq8Pdk8wPW0Msf9d6dH3hm/9iD5OQunMo8OqwxVQ3nHuYrC4WvelWOC8b8lSydk2yE/KQjc35
ql3mg9Aj3kRqT+qt/NHABaG/eP7bF0YJQlIuafkZTHS4X9CQOaewx0dNJiNeM3fj87cV+aiFOl+D
/elquDC08QbgIwrYrnI89u5jM57tKnfk9hIX0zqkQC+Md9tjUiEojpN7WUa3zC6WMmRN+6K6B5Ct
denZTI3+vfGCrDkiEtLNnJm2zWMUBwAj46N+hNDxu8weMpCUA6RSZBnO6N80rK0NZRJikkJ6rCTb
EgMo8r+7mqO9lOWDz27iA/asjtrdI84MXRe0F1zSLnQuhfXe5NVl5J3JKD1WxCq43ov/3u6QkHla
v2pT4cf1Cm99PxeEmWJwANTDLlAvPFSUe308VgP1eGaBaqaO8p7KAZARenWP4j6M3aaVWPv7iO//
uUkzYkaJvfnSeh/44kmKOXcXV1z+vsSVTVRMllatTMwWPD46XTXCh32wE51YOjjbfCtKsurlKTlQ
qR5qCxlKrxIuM00wszIbfFAywEctuMwnDkVuTN8p15DH07OpgNEXw0tWYK+LAgqlQL5kwtojSdm4
+Dw9aG4Fcp5ZRNd+ZKU1IVayy+2QYWuadIcHqymRToJQ6U2O58WdXAS5y8IWkXWZpRTbxLpJ8bNq
aia196CtS2e3WejQok+84apXLiXPR22WYTfYhhijNCU1GHQypjAjNK0jieOE8LYrg7Go1jXc4Yt0
+TLu2fd2JMHH3HUU+gcozqatuIfUPiYHXs2eop16Mqyuu5Kq4pDG6lCFAHOE+fFkngJyBA89/8GU
byav89fRZ9ckyARTzmszX8XLcr5ksS4aBQZGJt6p7BzcexoeQpOBMiXHVvHSbWZ1Zl9xOAOnxY6G
HjI2gswzqXcLHmXZC4H3D8KGv5dP958cx3h+3Ecwph/ZAnpandGipJhoDbxhV+IDfc85QyuCn0pL
lLe92gyT7Jr2SWzZwzlRn3nEfzhyLWRjvz7vubNT0XXW9/Sfble+cg5tze8UQYXcFczn3+4KTj1X
DiXoRqyKBjgxqlZ9Ek1buTQ23QfH+olRFGETVhgv0yAWmerd/5ZlIzRAZPq20BdfIIlEf1+8vv0u
aqJYsvxjOsIsBhPFWuQDMMiS5XncOudk6IvoRDuXPL+TQApzuwpsIJBMoqSwPqMTO7NqgusB+Ixf
eF8NtBubUj+/B1PffJpIENkAEVPk093Tiqa89d5H/LXN31C59+7usrlGrH1ENH/42F4oACP4skxK
hIm80g2FxCsp4oF+y15nrI9536VeEyTZ7gSNfXf32Kr/yvJlyWwpdHfYYffXp+UbWXXXFYCi+ZqV
D35+17syJJuZbT+aLEN6ArZgHI4fosRS4SGAABT75aBWzqy/kjwLONUlBjlBQbsj7KFkMZ8pN9Th
bBhAG9/Wbnt35ggwTTFUHw+ZC8nvO2gL6z9NIYFVSZrLgPK6LWOG8hV25kz736ur5/RbHjQf32U2
Hh+82HxNeX0pkZpSPnyo7qd3MtAmwIYgfTdE7/NwgYowPILRoBbJa/GHW19EAmM4Efv5F12xt/da
MkdDfBy6yR4DG4ptUyvV+iNL/R1Wd7Iz/sceLawjLLZ50xGDqpa4H7OFl+H87m48QjPtTVxyBM8p
F4ttFbLPMuAEkTI8TxgLVKNYSJ5YTGJzicxqa3JAY5DI8pKLSMBEMa3z++E6061173/qnK16V/FC
eV5BcZDplPJCwdjJB+68C2Ptu7MMiQ4g0ZmxT+30KWBfcONc3TmVZja3vffglNF/GSHXaU8fXRnk
XY+h6okO+/LnOb5JKevUjThbFgrpCFBNVQH/4QGWHaYc+StGNOfJpc+CyldVQWRgnvxAqdlz7+eF
lXYYQhwxDl0uizfiZDfLUapUIu84BY55rOrYU3yNOoSHbCqaxGtKQvQJMmusNQ0/d5KySJaeEbGh
y1RDls92MeEVP2HhJgYwOTFcU1IFZ4sOMtIVOAufgJdTyBFf62mIh2+Vne6aWzP/lhRNND9ossMs
HKGTaORw/ROokQeKhvOR6s+ur2gOgtpCV9L5cdQ7gGytYdq+lUSZbnW/HRZAaCsUG+5qe78pdEk1
THOy4nhNroAphIQbuPm1Ju2BhVjHIgnhe5h5jCYj2qe5z4uzr24xXbLQDKyhr6SQU6H0h5/VBNZR
xfyGV/Xko9fKzx+m1VqKuZ9roOZuo3A7xYafvdpP0cAR6vSuvlQWJopyHL0BB66dQAu8b0Wr5lyW
VRDpdyaYNEMIeCvErjPtdxGBT2LtR6uYPv83Jf9UKgS4AGUt1NwI2sI3Ua4zIAm2+wqgQXOcWEQq
v+5wHbry2+uOxgbYwEMkV1hWmaqecsBWfVmG1DFKYCwAhqqIdLFSX4AVHks9zCwqUJXiiHQR0Fas
prpU5EEl4uzUwIoC1/6lPtxCI2VIGpzuIcTC+CDgM497cr1YpfbLQvocOr1Lnh20VEv+osTPAk/g
l3MC1QPP2tBMKMKlzpHSKGS7ym+nD3Ms+HG1ke1VolHN36qZJBq39zmmHtEcM8eUWCqOkgQbnWdR
nqs4Qk99nDDYxaYNREtuPXLQepB0S4EbLOpJc8EAAlsUvXEpt4AE5+ldB9HmDBY/wIl0tLcsEN2f
oyfitkXb5Y0D3WM7tYFy3QVQqq1qsq2l/XJ41t6tELSNCr9AqXzryDpVwTVs7EBO+8OJONY+NFb1
U0KM9SJ/0Zid6yervsEIzsVtobqhNoqsGH8syn7opv0ebttZaaYEFXhGDk7pibSf0GxfrmCdZgb3
sgHMYe6QXosjRJSD9UHlurB+HI3DGLE8vE5NcDfcgLkORG1FQHKA/pWleyTAGMq1+VHRSKNxslds
SCRjREyMb91mS/yofqbDwbX0AaAbR7k2PJs6oqjEdJASw/tqpiOo9c95oxHKP2QaADw6hhFe/lw4
8yDmZTZBMjDOigVrNA4E6aWL9CiQZrGBA7la2RE2Air8oyqLPaqm0p9HUr3eBMJFO6++ijVFsmB9
ZGjQVcSeb3RCt0QhJ4RELReza3Yaxr/ZEv0CN2FCEi/gPBcuDBAbEs85ZV+WhFxHg2HyukIV+K8V
jtqBmlL0/18ZmgEYl+0tn6jII40gAUTiZxcCVP+1J555NE1fGeb9Ny1mxVc0J5mPCUiTWxhACt9W
dxoZ4Nxkt52EfLHPha7obJqtTvBCMxvwXPObme+014EnzSdVlq6gQLhP3R0oz4ftcf3l27DLf4qb
xmnnj1tm9SSGdhOqTCsIW5RoLYpoSc7gFAR1Ag2Hnj1tmzdAZbspGdMhNIqqyXgTPNEZ5736/Idh
km4mBdDt44rCxAaoOkhgvovAX8vIK+u4hVzsdbubtOVTqmC8KarSlyZ/WQhy8me+oIUI0Bd/aUgg
nVtLRLOA/Osd7sV7CxUz0fqWQK0IqbeHpRgggSRWbExfB/x202ZjGoe+jP97a8wgHMz21g2v/IUR
ItcWqNodyLtl8OCWiUsIs9R9koAEZkdKJClotDN8yijJ7+1ngxynPOXSYOuvLVVmHJl/a6OGIa2c
TuK9uo7b4mfVfoUxH/k7VkCi4OHfCvnRH+mn+JvZ9Z4KK+xLQbiR74k8x8E+9uk6vfscab2z79H7
ZoPzlF0c5dTZjr6vEVB5365YX3toLIUOIq6C/YvLgs43XCMJjRc/8rggURDnqgY13tdwK84AS9hE
tsJHcIZCSO+q9znGpIWsrsVQ6pfPS/i3tEUyT4kH4zBSEV9sAlAwPbvIDNl+7HvW7rv5hvsprWFA
4IJ0P0OPZ1lT8d70RLdtVxe/8ubiYPZugWAKCm6L8zRup3EVFXmjK0gYtFnLrZTFJaPzX//65j/p
UTjvziqPJnSiZ31fdbn2Y6JrsKL3xj1yKaBGHqV2L/P0rhisuagWETAPXNv0NOvlbfDgnWlnXjQQ
Qf67OveEeHPdus6cmQUUH40CC3QC0omIOK3UNRtUq4mth7vkwPHfRmOOyCn0QyfsQuwxYTTK8Ioj
u1UD3mLYKLJJJ3mgK3FfAokvkmzvD2TM1YNhDThxDmTXkPdeTeT4vh5F4J0XjbqG9O8pi4bPeKKm
ZTrzeAXjxSqM/LrcP3FN/NDhGY+WHmJaNQX9HDNbHu3H+CkZYG2lHDpt9PJQ5VSjHbemtQlI78Pb
JnkFQgeo2VGfXH6VNdO3XfipeIVm7s2308UbmcpmN6s38MiQDVW0b7jbWvAiEeWYnqkkwq15asKb
12T+Ce6gQFZleOGihuvPiZgvr09LQZ1dO84hgwE9Uc4aGtkXWJS1C4dpoiyZ7f+oh2Z4eObaITIJ
hjtjry7x3mgovX5YqYk259BJBrfy7v+t+LUDATrLa80ltRGwCR3dGPl0j+ObhoEWRotYy6YT54Eb
VRjqsVDdW8pDsWJOV3ypioq4NyQAXR8JBjose6UvOIH3Cpf1QQhT+1HHaA/swgR+WvqhjIr6rpU5
U6f7pH997zTTg/mAXKTZk9/TaDnhBNNrd/3yvR3jiR4RInRhDGr4Cr9m40tIe821nBwraqka4bt+
ARpkFMSxLJvpPifSY9oJ5xTCF+ycSldt5J3Sy7luyKvnCaqxo4YjsVqMn/XdvPNNszIDPgwSIwv4
JtwbkhMK3x8LhN2lv4d/4TQ2TcRcqfZTV3B/CfJhmnnCyzuQl+ha9JdL/hgNkESL98nxqa0hgG1H
Cdub+8i69mOOrFrq/sGuRp0aLLjqr8TBNKRrGjzMKx2Ulu4pmJokIzVOQ63xNVmoEVNY4tvTZ3dg
g8WEW7f8B+6dpL+bSHq+Fx2b2goqINSB4ef9HpUPP+hy7Wk1RzsGj3Rhsn4YMRRGL1sE5jfybtjl
IN8emZeDQQDj4Q80QyUIXqf3BJEsFutd2rv7Mk020wKxh1iNcQ24+fWCKdx37YEzK8ry2sOpiniH
fPBLX0NDkJkITEMZFezPXEg7cTnP9Rb60jHHwOWa+jOShsryAqquPN/7v65VrndENOUMuib1HkfH
0i5y7BCZIPshp57VNyfrj/8jL+MiqWSg/rmHO7UvzZ2gL7bNSzFvUc86P+H+cviXapTXms3d0v8Y
PDDC9fh+m40reXiG2GAOyFpOfzWlUD7h7+Ji8uBVE/z8NcgTGxcEq1D3qtmkQ3/w1kygpkZSlI5s
uyIygCwG0SzBS+7xT8EihPfDZtSdjMxbUBSQL0y3Fe9MRIu/xvG2RZbr0YxXUmJ7CHg4khklpa/b
MH1OtDl3HEKiXsaGuoe0chbx3jPRPO0OagVNTjEo0mGQw/n82dFC4BdbJ5+pN7mVe89sYaYipDSr
IZjqveCPDLJGdI9y4FwsscRSvDizq5nNYR4oVsBzDGOMoGi5yImbrf0WOBvOw5a+gcYOZMgv2spF
WNRD/uccWDjWHbxix/X7HQXHU0EuWnHwLAQlPIUwo8UTVrIgumPsjgt8nb3An3faSfMwrYZMf7yZ
6Uo69HLDwj0FA5f3B+upAN6F+kpQFzKZGu4paf5nZu1osccpAUQBkMm4S4oxbxuw3pHTt2YrswXy
/0OSxut5CFNzcbxqvHOGVN9rgQ0VMurKtC1J0fTs5fW+IPDmPbPiqga0kcd+0w4Hpu9HpTbDd/2X
RDU/RGLl3O5xTbNv5a9vCF44fKR7FPRkXnswzdwz9hO4/uN35M3wjPUfpFXGM6ol9fRnnuKL8Z3j
+L9EcaqN9mNvAtg1Skbg/YKPg2NSTcz7rUWqgopBvslo5n8Nztpv2aSi4UzZkSPZvHA8alyjKYGs
O8L0ClvQJjJX5X+N5ASw6WN6hX0lXAivj0/A/Pe5F79CO2/A22H/51YyBhMpXVYu35KMoGdVyGwp
8CxaCyP6kAVumustZaA4I2L/2Yme91q1XqB7U7ZEGIKbxqUwvwkMb78y0cxHkSzOskUNUvrtLXw4
L/DmZJWqo4Pqu18vNtWJPJwj16tiH5jS/8vBL8zskzhHGbppBM+KU/xQdu8s3F6l+5o7hm2sTWy+
T05Mbe9vhVGVtVK7Qw04U5H8iPgg2OWHFI9U3gcC2UBhlqXxaiUnATBKB4UDI5iaoZvc1YWyeo+r
vbZ3ADvCStrP8RWjuCTE6VIUmOP0c3fVQkMdqjF1icbS7i45dinTD2DEoC979L9Ry2HKQxX62PRc
viA+0vv9GEihexKzSlrHpvwixxKI+8jqQT8dUvfV533nH6uWzyBl+0R3OIe8dZJTnxHnalO3mLL+
jwwaRuGXEcLFWgo1aKWuug+UvxgMGWnE3Jp8rVLmFbY3FqpwVuhKVJY3fxHiv5YjFSo4q+EnPk5L
rxuxrLYk7hg1oCXKEIpaEUIkjySL/l+i8HQTz8nP8wMVHvq/ApAhg4Fv1hJhopVrZk6/f1j1bEhG
hjGM66r2dPKDtyr5Hf8zQmq4/QWABYLIaP4pVuFgH35AKR0G6PtNmK0XYra5C/9+heLAaZmoCp6w
dxo7ujWwsZ+a5moePsXHhxsPOBkcmaw4Ce5C6OvThkkThYvexkwKekeQMs3NIqItKfu9OW0CC1eM
UEixD97d6RL7KXvOubqnSzNb0X2cTTqBsUz9Ps/XujDHvtvWWSoax/HCc5XAkHUV58oRq904XmKn
acRJmobkzZlm1m6y/XhbJ61nAhfExxw0kB6zjjWda9AdbdiP1zq0TWAg+MHJhAmAGI490ZcuCLtd
VRT6Ym86KBOS1aMaZvgGDFNeIdSpodhQQrd9PtTpEdFKrzhfSKFcsI5e1DeWnrEKb5ZzwzaBKEGf
sr8N13zWbTFGAPU+301jB+2IZNgnLTIkRY2ook82rly9nLvKb0KspmfWCM9MYr51J4nKjmWYWzL1
sech7BSSzvI0oZaJkJ24qHwTWj+6rO20ZfVHZEgxrD5Ci9VdC8xrSVZ8m0wQFVgTYSTq88s47lJ/
NbinIEY+e31WHOG/xRx/okCuJWZ5jHubbI9Mi7lgrwPJb4D5ncCYryvyRrXBdtvHKR6AiaMkv5qw
bg3NujBEluik6tvWYl9xxo83GhAEXiQVkaM5F5Z1hKKHILi7UT5L+dPUukdCFfmmF2+2C3auvDgw
Ew/e1QNxLJSt/wFVdyWlbD0PtBiz1ugnnQOanQJX4LKs85rf2urbvAeZ/nkSRIe9ZBDPkRoYXaMy
AK7n3U72Jkh2dISrVK6IQIuUF3q6lrRprOmuIMO3iE3z+mcuau9c1SLg8Q5xtdC0qmQ1kb/HXHwu
K9mYxtNQo/JGgiccwoQ6Km3Z1f6IQ8B9ZoEwBrj1/CQaCnkcJ6aNiEd4/lsPX3FxS7pxaJFyqxGb
12mVQ4lcUMtkSoH2wEUURUlz+JiAM+Y1bUJpuOjba2ml2Gtjc/6LHlFHCPpOtly5YFgTD2SmpNPv
GHG/GIZjv0CR0gUShfVvn6NqpasTYkiohHy99pCaIw0+nZ+iSzG6fi0xZ/vAZI0cb18MYZDFb/eH
l+IyX6Iin2dMnmwGkDvDh2SbPlLZXKiyFnZ5V6gwQDRll1C7JJl0VjA66IP4ne/8h6PVn4r+y8hf
spALzIim9Khrn0ZuX41fQDZMteh9h2Ffq+1MxVNtOxfMpDI68Vt1DS//c78MCUc0+/Hg9LEWVUks
4qM1/wHPTCK/QUw296pER32yvoJFGhVVMG3N+9WRVg0q+vDG3NEaz0CwhTEHssQMnoGKD8b/wYTN
9zdYy20VxKRIb4PY4RlcZ5xDMCetn4yDnfiSlmHShPcw5xOicKFbsRNkN3jAAESYLxbd7gUs8Njv
nCQbMIdi9JKdHojFAOa+x59S6uPcCYM4HV9kYlsqWdQ291WsyTqOB1EGEp00k2pD9f+PPmS5C/5y
7bmF/aK5CoMSyVxIQ7OTnXblPGW5pwqM6WCrWEOCT31CeLJpf8sMnn9WhDCziUcC0qFrXVPF5y5n
5koEYMVOncM28BFO1bdnJFjvUFGsKE5bK3tNbWfmQYGvzP8EvEDyVS4kE8ByR04u22AcrvrZMH7w
DeSF0b9x3sbjQt/8pxWAbCzTmKY5ndJCcFStIvBNetpzv11pFoakM6zS4Blfxyex3Id5Apl5G7b+
hAnctSSKrmQKLdRmsbqjoFqJ6Brt3mmulpG+4kVSTCxKQXuG+UxpdSJ91h8rI2MZ13PrCOQ1BKjh
1XleqnwVeC0It8cCZYSlVY8lTPXUu6orilOTMMtIGgn9QCqLlhceo+UXRKBq+S38ZBEpFbW5lky0
MbLkjBUuX1g2TqnP1vFSIn/for/t08HEvETnRnn/o6t4RXMa+1IZunowL1JKipmJQC1Igk8MPZ4I
yjqPhF7Rn2AO2F48gF9MqL7YNjLo47tX1Gj+bud51K4fF0JSbm0mRBsTaxu0dT2d33LFxcx5vSDd
YxRW3rGfO5QVzUdY1bjSdLFMBLUVgNjQs8MUb5SFWDWnAXFoAw4al3XCY1Y5cRtgGzzg3+MR2Tjk
58Qcu6/UFnfU3m+YE3lZhujdWSgxzetE0m6hO+5Gumyvk6TK2K/WTV6YkpaqVIXE/HqaOzCDTDeP
wjmGA+R83QymKVbga/639Jd3RBwT6JmB98AgTbTIz1cd3ynprW0mrXQMebS61ZXNzWRXHz1gmxzI
AF/a2b08/FYLMBrKPWNev0i4LyKsvkpCztcFU3XSLCWtypM+hJP8ybIC+1CBrBzBS7+DE+m6mv2h
V+kRLOW0JhK6CyGR2Gbbgu/a6LmLKEo74vYtXbNUJ/Mxu+jRKBc/pJdLNeOxcyErfI+5ktqZIiKj
st+CWyfc5UDFpbol90uxUoO25NSmFmi8GsAKYSUQDxS40e+YZONCjW720GweOqNQbftl2sAy7fFO
xu+pHWfq67uMT24QjNr+FejFDB2gDrWkQ+WwPHrPo7o/jBxBxUumFSVrinwT/TETMYlCNrZNdx6j
t5hAS2kVN4AKZSwktDpzCkZA1m+CX0f9qaw8aRreTthf2Mca6XmHpNXHUPL10Q/hTtTdgNypBCtP
plhBUYN5WVdXwNIkwE+3N24z1e4kAmuOs2It1YPnj48vInCiF3gDo+HXI5gnSweJzpLUHu87H0Z6
AqGDjXa72rFTLAuiBo4RT6CdpXYCe39EmxYuULci/u85JhompO8ouq0ljk0/q/9FJu6WFL3wy0le
tU+rW7YKUCfYmdIzm+f9WCp5VI+5lo/+Gb0pt1lBTA6HAYLdCUNj+OEv+RFPiMuaX9BNHMhREbSJ
Cxqjobay9siRxEezs6Lp36QFoRZWYyDR0iJ/gdbz9TVUoO40NPlEmUzALcbJvZNCS8O7eUCzMOZ/
KZYbtTjplxhA7Eu3YCXvMRNYaMWdW/n7Fsc6UlaOj32HzRpzx0ndd0mWnzJ+IOa6LZENfsLq8gQD
0DMrKAQn35VkMTTjyrHMo1HEyqcpuIWsiXzDm5A0bXdiJadgoLs2zXI+AdEDW0kQ/d+XwoOuW2Dv
yE3S3VQQJUHvIg1vbbYsqX+2CshxzKwKd15dDWjBynIWIiiVMhmJFxxfs3W3812V1W/Gua+OI5SN
tpfPxLAezNXoRsLWMaXBJRZOmH01bFqAqF6HkzTMUH9If/ysMuF07ZYIyeyP0OZtRubcxuBCFSIm
3qubtAakJI1NARb+mvAZ7bBYUcDjjzVcnha2QCHwvQmdR3bfRFqBnlvQn9M8Jv1nT3XW9KAZWV44
um60eew0s6qKZ58YBOXyh57nuvOJmVeqH4mP4Qw3vtPKWWGX1SvC1lrGtDZJ7j3IHc1bSepQeacd
GAyWDaFbwxS7NEGnutvFxWZBwYe/scjIcEDz2WvoupyrMNsxNzpWQI6Zb+vIbFdTUjNsz8X0RlER
LOn03PAPyXLVtuyOEBmzWD2einbbzT2bX27EQXRVqG0Y+xAqvTC5V/CcGFBXZDUzJLd5x8jttLw7
niQdNlO2DYPI5gJ7pq9JHyx+76f1wNri6mFGW3QprWBFCr0TpgqtxgWa/9K0Y+O+emO/HVpzrnlR
7JjsdhKpL/AYX3qyq64lrynIPMbVNy3OVEYeUvyHcIbk/6X+XIS1Hq7Scjz9Vf8FIYBSUl9Gp45Z
VPIdBrfo/x8rs2Uair72uLgYxfV51Pq9zJMVxfsPLiLP0chOZNHMonWxu/lB6rYKPjAF8vJgC0jE
2pGu+9jXfNkDTgfZVKj0ipK5lDdOEm/GcPB5yJmJ9CtzYFsWG0flDLlVqRjfbdH1EPoNadTYprDg
jhLoMQlZmBl33itsViH8EtTH3oYeGcQEfQLwr+qbHC5pCNruuCoGEPUOcjYSsQQ+B46VH7CcSt5e
8MdHBdJ66JflOmlykp3ooBBLdysST/dP/IVB4eRM7DDk+ACNC+KejiX7kfUM2AeCDA/OCfvjjMPu
qLBC3OGscA2wR0EIfpAA5kZ7MNkcxSP5tJlcBG63Bi547Q7/Eb0v8/vxeXYt01MtB1mkpyTTuBSb
EMn2qn9lHG62slmcoJo5vBAL2XJsfPuitwKL5xfOWkv2L5eSaB/XpmBXxaPbckB2m088AVTOZTQu
Oqe0r7ViNg/Yq3sCa4VsolMh2Tl135rMjLJS/yJjcmPVt82x1ZA8lE4BQsKhUwxhYYLnbicJFFj8
KRkWbUPxiZBysi4D3wYmHOZAIzJfhOaHjrSH4d/bw529HBjDZsxmN8hm+4bhrgEs0XrbrGfk3mnP
WfYQYxv9HGeAlo9bpsv/nTsMztRWtIA2RMTkz9QswSbpZG9k/4XxTaIJRpWC+K5aW67dwiimfh+m
Dq82ybK9Nwrcm9isum38FNd6dKTkE/WgNGJzk7vtO/pQSPRZjmWXPmxS27L097oZxxrXt6hBiBM2
MaI8NxmL45JJ+eOPMM1Rot1ZUFR7CyYQErlytTpZdxQznM2zc3VsanxdABfwy+814wailn6QRxHf
QJfxFWfPMw820LBbVbHLafRYJITB00I+vI4BT/uhFlwPmRy11I7e63jb2o7+SHUcpUUaMNmkKYIx
r+Wjddc4tYXwB5bCu6Y6pu2IM9XiLi8DFA4fWH6vrNjlYG+ggmS+MHMghLWkIzmCeQtgv1+Rennv
thFMSz5v8rpZ5p7J/oPStkLD0hYL+XYJYUrJUSMkaHoTy4THTiFtQtZ5oaq6sqoABHRdO4EO4YHd
nAkf/zCFhSUR6dJWJKaX1Kj1dt4Aq96vGgMhTRaADQFfRUqZuXvxTRk1a1HgrNxWpdGLqnKamSkc
xpTBar0z/kc+8ONS3E2Ge0U0SNgovgdJw83xyZPg44QUMU5VmucdNFHrtDrfJdhf5cZdJbwzoUTJ
JhaScPNlrqTJjgLP3wHl2MX5vbPvkqg/im/G/nVDLU+WjKPjqAnmmg6sm2dilvhrc42VH6BqfEky
5u8XJBZONvitDmIBNqr6s8oRAkxadqma8c5fNrdwU6in8WupZ7S4TXQCyU+7Z6P4c0gOylpoVD4u
n1Jthnp+7ILU6KitYWA3zCdFRHxqD+9y5Mj2mNL6pn2nfQhuLYwaHHpYCSGeZw913IzziaPFeOPJ
ugwAOn0TnKiXSwaHIHWljeO5zYtJvaNlQAnpmOIOu9okiM3GlAVMfLzYq1c4/EXKp/wt86F7WPPC
6V+qC1eeRRlIGFnaUFyslybU+hYdOC58GtvKJeXq3khR/aB9ver3OGY3+JCNK4QzMdduuiEXHpO7
bNMPCIjPEGf+xIswQbo9Jta1lQB0jNXkihC2HSqsOu2oS7jIVNV9/ftzezBmn9QLIqZDJ2FeCBCc
DVDL7DLwqdyWK6eFyUv7a/a7IqPK2Cgg4NsWEyJ7j58kRF+vThFGzKUA/KxoI7ZezzzgsWh9T8x+
QKLeCj7bFtmfKXBpKNg7LG2tAhS161PTFbBXv80sXPR42vyP3uoGHBv4fYWGs99Mp4PZauGII3/f
FNKPLNJrXvbwxVqE+9ANxBuEpEqHTY9ubsSzaCKKLX9JiPAm9kIxwgctJFXacMNswBuCbn7v73ll
pnePUBk34qT0pz1Hz8vI9H4z8Cak2BNilt5lwhh6ecfkN1skPB3U5Q3ntU5CYw1Brc2kpPX23kY+
yJo7sQ0FEmdV3LsafbgiXzjT4WKlwq77/MSmsXqeJiRL+hyQfNp06FIUGwMP0ypoZ+ce4gtMj5W1
hsJugzMz8cSBhAvYq3m/TUm2oQS4sf4Ia+7B/Hf8uq05Pba1SZxmvH4zyioABYqqgmOe7yuh955R
Q5aq9ZZsnLHCE03NdymgiFUe1BORgw7yEscqIdCnf9oUKOW0V/jrpzHNQ/7+qVUqiootZrQzNOiu
d6uXfPMKp5xTe71pa35RjRWqXjVc40wDPNeQibzxzwvuM649KyZWJP/di5pIqANTX7LIQ38MScBh
3By7K0VLx8oElkQqEN8S51JWpdaPOXXU+bnr+KRKbO6qKJWecmst6OBDPevZ+Up3jMLHWg7DuKML
Qcj0w+qP5HH6bdkEwDcW4ijyd+kvIiNObgOgssZEq6sBYQ7PJlAT64motkHQ/myYDVOgi/JWBuO+
oLGM/BhhH7OjGU1clhmcQJXas8swZ9FMP9/xSp0cQM8UzkRQXTaPX/IiyHWyZ2i5AwyMiUW4tgLM
hjdKCkxYuH3ST5mF15gX148NolhcRCdQMvrqbTA+S+8ASKMatlWDaqss6qRyDXuWtyvtYQmgtpt3
0Dn9iVx1Ln6LmGgpuTOxw/XVLmIuqSCuUjSONqc2QOEdHHlHeLaLARMa7lqQUjsgHkDmNbh8nI6B
Qak4EN+9yOuTrA0FeXHv9gCyTGbkzathrZ6QopsR0omKgFzHan+6U6esIpXaLfdfkolXhaEY63Sh
E3hhJl33Sng9IJiFmcaNIMJW2KB19n81VUwsxzhFCHefaIcM0WOc7OR8nSaqYPdlZ8hfXNw4d/K3
SrfOvI0D7obv3AyZX4X6EdrOfiUrERVn77+t0CTTmVoHMzbA9BYGl80jRy52tLW38bM/Kv/Pg8gV
gPzJUa7HaiZ3yOOHm+Ou4WPbQj+NsvAoOzFSUx1jNvHwBplMvoJkRoVpnuovo0g87gCsyQpU/5VU
0w+No/ibJbGmO1Mz4mjEUq5AGy1LZK6D7t6EY05tr1F6BIHyKkcjAb8o4FczpMyn623abJiobptg
MbaaHfJWdEo5Tqc1PPoyT8BgqY2r5wa/MamZ3kYLm7h4O+l+qCKPA6M9HKCWOqC1lSCmWUGNC4ao
zEyN8T6ZCbhzqvTVF7ZAAc3DSEoUoXPzQqX1/FD8Q4alNkxluRd4COMlU0jYsC6xcsHMFgdDSzcK
2zApNR2JzWyOmdRcoStrCCu/lRYMm/yOdi3Yd5NLD8IjtjtnoOOBSg3N6sy0/cZMHe/qd0kG/y7i
DYGTOcUijfuluCKLUTTaasRiDlbPivi+8Ag3LYf61eKoAkud09ZlkadbM+gvoxNCdbd64USLoGme
nzbY79lC/fUkfycl8b48Zt9azN0QlvIqKQhKpmasuQ+dbfxhRciUtr7lG9eIovfLOik9KyIceuiA
4jxTkssG1DwCQU/J45ydGNfPZOHyg1ftls3vV/DALKKFCW9M7y8A83jSvq0pZgMhclWAwFHK8TDp
ftwHD0OR9zz2qOZCXLeiV9+5ZY7cnG6x/r6i6Ax+iMQS6F+/J+NRpyUyZ8ryQ1612R6QxJ3Lvci1
MBl5TL/G4tcUhivPmedWWb0NAmj4vtYR8DT1Fae6Mg5BPJ9N+ZuQDTAhKLpFkqILiIWn49FoQGF6
IsfwEBvCh+OvFWApW5ROF/R4YgEdcccP5jiiodb7F8C6h+0o4N8zERboAhLT90Ih9VO/yZSbV+B9
Eq5qyxwDQZfWZsBYmG1hyEQKv07SegZ9n6sGAlp2oiRTC0RgY2m73XYxzVurF0WK0lhgHkHHjtth
kD+XnWmkomu/1q6mzFoCbKDDXniYHkfyy+A04an9Vm4gDKgwtZAHg93I0nSN6rH31ZzAdfcUzZws
TQQZG9e3geuMUMJ/sCC7PiqWLSNL/+qq/y2+BAcNNlp2wS2XbYsitgtPc+5NQtZUb/uSrmyqBZ1R
u7liXfYrjPgZoK7itbV7xPxoYRvhjxd09X9pOb8epH6DJd536LbTIoxa4Wnq+wSuKINgjYOMJlYv
/TYwNj6RqWjS7NPvhXAIpaWzZmgdswWIPoIg+2w+rEVemGYu5o8WsZFJ8A6+H/LWyUGBBBlBAkgy
BZVllOJyLy8O/ZcqKEqFiIEPbJMzdraxQmjDefmOK8UBEyq915n5BrftnOF88PVjzWoXi0R0bJ7W
Oe4m/+KkpLlFsvuR9ITzmrPf7ZUaGTmlKqRRoOvm/Tj/tl4FLIWt50L6H/NFL8eoGYlfgiRDltQc
pdAnjAfbi6aY02RpHAqXDcExQEg8NoVFqjvl+ybqs0Pu908JOdnp7FU2slaiDqaZC3LdnukMGYRd
3Z5VES2+ywmqdKrsmlJJwQ36zRWLNdXZs/HKZmyycAzEdt/77izuP21U/XU/apW/mSa4fovSPsU0
Vnh/LkUMfwWiUf1+7uBOtaDpOYO+ZWtnSSr9ZNELAd54F/HDu6UV9DhV5mBAbG5COfWJQ9JQY+du
JM0mjQg4I37R3ClBKijUpzDtTISYol5LVPVMEcraDM4N34f3dIxMH9dcvg+alIGxQ5/nZcFlREeY
2DQUklB0mNz04TEL1NodY9YDSISD+Ey2LA7gcxGyaTkXlP6nVYBRnv3bgL3mAHsbbEgrDxJDuNNw
A53Vk1GGhReFce1JtPUARUn2SdYhVDBMO+A7nMr0M7TkslkqhdtDzIACo69gq1R4+6G+6OJrotyJ
VqVslNR7P39nX9iHLhguQha/fS96qeBvdCKO6gAN3XFw7RL0vQYsHhcnGaohvCUU4P05j6rJS16L
QHSC6VHglx0Vkw23iXRM7x/qKYtIzwpQKt/FomSJ6zk0AnKDd1dcKEG+fPXQKGLv27BbhBM9N+kn
rDuvcEePpzLttlwfO2oa7F47EbadBhXISH3BSWcKFBlQfmyZy0BPrx/+Okb7OxRu2DP/UcfRNHji
P1OhzJlQDvuThyOFq5Q93iRf13d3+MlpBBLSsCxGgO0AhGze7faAriQhE1kFeTElNbnKa82qoj2F
B26aTCEWiMhrHpfSo9UFaOaGLy+5MO5pG4DQ74uwguED2INp5I+5iELpfHDRPMF9gWtRuQ1SPGlN
3fRBXcLOBWsG+Ytki9ce+iwNv8NR7MUGztQVCqL/Ij0jpiJMdrx8XaaaigJe89sUwFTZm5L4wgL5
PiE5cB3Xx3f4zTHNKdYgZOA40IGejBWu4IesiW1zEVX8lAJRy8ufQzCyRTlKKiT4SVMTR9jOkdPm
8HVQbg3FRWS5s55GZU4pCmnDn2pN33VIp6mOnNH0nvmm6bm/swdsr+sm20EOGjBGLaCcjxlePIDA
QmTkRo4jtdXHnJCWBOiOaKvW/6jF32tpa7HYnNp+sqTFXqPClKvo5H3iVSUArK1xXBANHD+zRGCG
UoS+ivKYcHKIFiLvTPy6z902F/4auLuShsUIC4Sf16M3g9lL4S7+X6TTSY/TSVh46kpqhnwklC7g
vF6DFMZEcPnPmVog0zB7Xc6b366h7bQwF0H1jm53lVv/xzaeW0l6pG35BLt+oIQeqNjCtoNOfoNf
aKOca+VvDp3DX2QPTam+zVCd7QksVvFA9rdHTrRlvInUJrDXOgWnFzSsjkDITGZDAz2ryIn5NSTr
FfoKS2ynSvKUcecLPqOClwmRypvO48VPtQBfpvxMcmK0ggJKxPT9+rIn3omPuS863E0/WRvZtULN
xfydIJGiG+K15t6v7oqdUm9wY7bIbBh9OuFh89umwtS2QV5rD5f1lPTKdKcmjBvYxXoAt9oSb7eV
W5xC3IsS7IAqpXG6NCwFtTHhj/vT53DpInnwlfhTSNChqdGATpK2M1U5oXpV/wODTiuguHvQDVVx
wsg5fapV4hfGwni8+p/Hx2bT2Zt/QCPDCcyxT67emrN8nMlLh0gaRUD0h2pLCjQMCNfrPeCU+vWP
lS82uR9i42zKvUtg79BHUkxeqok8xOuI2+73uFB5BHUBgTm8+AkyPOmQeEqf3PqSIKt/Ui/iyAu9
um8lpR7flrq5mlclofArHfdVy9d7k8iv4CuunT5EN9ACHBsJI2fIzjOGP3n7nJHybPcEPQa/2f9w
QcLktiIVWRDtYMeuPlZNV2H+dRoSGzdJ1pfrPwXg+XOt6rpE4BHSlClkR2a84jrfpKyPcbenGg5I
N+9I+ERbq6/9fjaluUDVbaaUqoBMDsuenelZQ/mPpahcG97IN3XnE/3yVKnZRSfr6YOOJ/Axo0nn
EVjHS+mTbw9H5tsHqx12jmlA4R2vyNTGpT54r1KZaZP5EeFNpgrw0EzF852iN44s7u2QBuy91eXw
6u+lzRkGZlyn2wLti1rY16X4Lm6cJiXdzZfnuv9JM8gQJAGUYaL6OfrbduND105sgW4Qyzxl64YC
KZiWurllylz9nQLImWLHYcQ2mtlN6mOnBYXVk5rni43IiT7Xf21lit/DNaumzM/l+7ebEVJR6+nm
0zmOZOI7LmjNROzfm2huYxFGdsYtu1h/NE7ejP6JMDfA346DDJgVJTBKYV0vKxB5/8mJjPuHfNn3
S0Vjbk82XE01HnimiNyPZ693gDZkrye+zgkLQlqkUvq2JdIDNXI6wwq0kp+vUoJCMzIoe/gNhEC6
+2Vm2dL6K+mmXL/ewCab78/JAfXbUmt9ioNn4Gevm4RZIkBwy4hipWNftc9wGp6aSXGkVipjAGvn
DnZo0t4GFVNqsQaheaev+TPvytaN24lP/A4oP7aCCFytj2mF/guTT+4APshBsnIgLGNtcMuU6hwq
1i0+hXEBEwgn6K8pmQf6F0zPhkzEc/QgJA3oSORMLNlFS4+wUu3V8pSUmnW0QgPZoy5jUl2amfSR
l/cBGxw0ck03Q+WEZi4ydzMw6brY+7PNO+qoYYxoSBiSSUQvAZhzFEcdfySDswgujRrRcM4uVjlW
c0Kt/reEEHl/1OdZJQ3IQVxBvGqlXTuXsvoyZL7QYeeJn/smocz+vsZVTCJ9YOQs8PGjt1zI0z+h
eiq4F9yIs3el6H1wtr3HenSyyfNeomeug0r5Ib47lQG3sD+nHP06Obn/84JKmI8rJjvnOwlYL1Ee
fUzF0pp/pHLDnBh0oRPqbI9aWK/UcLjBTnQCWFbeBjDjGU0VOv0a6V/sp/+CIw51mXsG+IwvuYLr
MA9Rd7BTnNMcTKTlSlloeRabumz1ja02VMeZ5IWjRkuocC8kQM99Wfg4y0VPv8ktkMFWRaqGDmXB
jzBJv01cDwAI7DkuGad8fKmz2aOGm+zmEPfj7GvqStXi/6irucqIPTX7prprNe+T7lNrTDCpwDpr
p2wfRdb57yhQdwxakZQeLqpP17HBrVN3sTqIChCdhRfk8w7rSWpTlPu0yMr7RRUsUZbt6uhVyaaK
bxCkDcQ1lTmGZCL3CEnXAzZa+eE/f49qbrRff6UgCVWJSefaDgCrHCTWTuDOdHEnKwiBHL2vtfqI
J5rC/UkltTZ3QzM5bABqf52PQdUurRDTjstX/6czSU1ffgVIzA9tFOgUmCpL4PfpAyodQmbuMGNq
RAMEcnpMvysKfixWraCiWqyFXxVd4fHpipJu967DqvjP7vnIFVGHhTLP57AyUMmKisYyrzepAKfN
zdTIoG12J15UuC8LVJPXC41WdlsjhDRxxvuMBY8lfqPY+bQ87CRqDAAtCDMD11hbwBS8C3mh1S74
mzB1IIisuEiEaNAC5L6FcJZqSK+dBFMpg2LF741HkD9BRx0x6bZlzniFjLF5qcSBqn3uZU84e4Iu
bll8xtv5ZSX6BcLX5xdNHm05NDX9Nv/OUSN2kQXm23awWyzKHFYk02yZEYw7wATZptH8GpdGWkfD
nU1AFm7LPn6cYU2HBzT5u0JotL4K6ZrFeEj6FLXmzoQ33Qsba2p5xay4BAUi04ndqMiSPMVcTyZ2
C0+WyMa4wO6xamA0wN+fnCBA0pAy9z5wrmQh6SJGVKqj8g9GnXGiZbeR5/ZWIPmGuTpnKy4ygOLI
o6+YSFEh8JGU9SIP/4K4O23jaF6DQPbFj9zRQd9iiBID5rVdtAGDWdyo048u82SSXFejN6I7y3T1
6aWdhyZVLW8YtfsZE2KY5rsyRjHh7q9vQRuc2aEkB8122cAGzXiyGCw33irBnNCNCdQnsWrXrAyK
P9bAkAZGKK2FZ8jy3ZY7GZLT3H6LECCFYyYecM0QsNiHzvd9feW6/k+m2qDmPfpUU/C27qsSv3jg
GpY2mjrL0M23nGhWirnbT2STD99JhlHPI/gtdnLg9L6vVQpSg/6N8eaew0tx9OWvEKt/aAchJDOR
DH9yrtZdnwlodm2ns8FPmX5yG0FBHr9md/16uSrUSGVw/3Sc+U0srhWGxSQ5VeiFuriHA2+Dr0Jq
ZZxLybdcHiI8gFsiPQs1LYCoQzt0N1ijsBBdbyBR5LvqQH23husRfyhgbFbeIWAwAJROuh6Nb2nA
M5/WCPxADLt4UchAmAcWxsAAZ8IXhgbUTmtbTK7xgwzgh0DgbSbt3Sm58g+KRmYkk+Ksn9cANx5x
kQzpaXdM4oJ6A8u05HpgSAshe4Gqx3umXrZEqMf3K7bAw05M4hhMTO/MWS8I2Lv/1qsJtHgxU52q
1mPX36tsoEepQfDrrKZNPq8XYreDQebvJ3b7zb8gXpbbiF3MY1wzppcUcWpAnw1FL1ZPtJqQDO1A
rFPCwBjf9uRsvVvaSmR5/nXjSNoN7vUb0qIzyOD8WAYYyFnL6aapRXZSVg4FsFTCsbESjOnkjee6
VNDP0szka57nPeoZ3daR5KRbyt4UAkuCwBduhxQZurHqKeIL93AtKC/ecAOx3/hnSOJp51pAGpBB
UkuEbRHQoEzbfvP9347Ko5YH1tlknBh6e+hHR4kdnUyzGnh1okPumfBKn6Z7q5MvtJHko0WRf349
5HOHI8LQcAfemxMwifC8GgW/L+WK9DPtB9VsWPalQ2PRKXsMHFwmm+fZhw9Qyj37AR1G2p9jmlM8
E2QNcw2o1WJMRRDfwUS4MjQWhiPbesmaJV0MYWAbLnDuNU8yH/BzFhejoyqU1SM29T+8lPAVwXed
jETFj0NVAlbJWomPVP+ybaI2a2ouTYh2pfoIy3mkINVdF3twn6PBLqdqG3RM+8H3pC5qJwcHL9tN
/PjOeNWriuGmFKQSdfDd1AKfGjfaW4oxpCmPIXpSD2lAxlK0J+hQ8RLxvYQRT8n0QbHphg2z1IAv
sWovtkFevGoqt/Csz4ukxpDJMPLsQT3ZocPAWhYezfhvQ28ELrsWy9px6Spmq2ZiyB0uoNWxWxps
yTYwFL1FzcU4y0kfovGEnEG6nwxTvrjpFN5EbGNy83/qMzFWQDVZdpS86N0+4Zo/HmwqDaNA9DzG
99MmZL1Nwh5CavE0eAGRO+jyGf0lzzS1BZPI2JCtOa6pOwfUEMzE3znCJRtmBJB6LOFQCdJ/+oat
WQBghVQv73sO3w7dXTBONfqzponBCIOu8Aith8fVh9AlMEz7sckYTNc7v9byAo6vCWUP8k1cjSgc
YgbPfiRUXGByG+J0HaKt2GNMowv/hvfwuJiFKiUy3knIh2TYe5nDF3ndAyCcwLplSGZ3i1URprlg
LKJWzWbHZRIeC1B5Wdk6FTF4XzAMWrQUU7enAZdd+ZzduHrp6RJ0moC8gzyyldQTP/sjSGuxOfvT
fmaRVpV3DGAKY72kM2JkbOfLgfNCP4+1iVV8Oh2rJvfl7KspxDbjyW8YZo3Fpv7Ht8RMseLVuIyR
fmuH63FP/A+COhlaR4rfedik9+NVY4+WRsVtXplPOUG6tZcpIpv+X/EUuH0E1IIv/XduM/1CmtBc
MqrEnCFiTDPQAxJb0/Zjp7gHBAo2Kv6nexp6Kqv9yqvkamXQN+JYdwIhWLK4InCV4vPs1ItcfDot
zJ2EETK3KDA+lUXK39qCqishoxlfRJ4pvgAvjUkeA+D51zg7H2DIEWB3VXf4fBTRgYRBseeBRAlh
xInZrLYH+p2Rspfijx/lvV0QozWjh/YrlWURgy01TatNF5C30yZaWqJIGShqmttqJRKoPkw/KNAP
PsCYW4uk2xxKJCkwbyCMYgnNqBCbS+Yismxc+prSwlHv2egib6dOloxoplcvzQEFOfRb1mddOV4K
nV2c/hXYDGfdWOkTVzDUnF94sy5QjfZVy+Dr2iz9R5czE1x6X81f5Y2sFVXWNmo1AAQ2pkMBtqbU
WnH0kDfI+RYuNeFepyEltZfZs9/Y9bJeHrmEmodLmhSwYQeCK9RKflvjXViSiXJjqtU5BOEkuqbT
jA3Zb5cYcsGKVmnk3/A+dZXl+BqTywMGTxax4ywhz3pRWgpz6tqrAhuLiHhFn6AYZeXuuaLITh/3
AT45sTJb+fYYJ8y7SjUoaEtrFQv7zxGA3QoS8NEejUKqjrCYw9VWtDdga9RHnSx98VBr2Rw9TOkI
JNjWsjyyGcBmKph6v1fWSgkMm2GI6fZuLDbqnhjW3Ei96CelBsGYStFD9+S4cuv3TWaeodYzbhK4
QfiRJhk5PkK14Y9uX7nGEL2R4x8vC1YYKThn/HhFkkGPgFMV9p7eTqvaf6W++FmXphmD9mQE2Ef6
l7B0fIm9wjTOH/UqYJX3f9YnL6jNbyGAi29vLoB+zc15SzmLybTnWRA26PgWliUHVcKU6tV7WIxA
JFK2hFZH3whwmqckUFhVpJ+8qdVg37vHxABEzMJwmn4LSbhoNDOZyCSk7xN7vCAy7HAFM0AmKeAS
DwVcfDrYtDj3oWyBtNyOxIw76Ln3WxuobtWiFC4cVLNaOl9tuZOzmU4WG00TqCrvZagldruySpj3
R7ja0Tf2YesEIaDhzUzluIiRI8Y1lT/SRJU7dY1bjgDbaQhOOBfSdkiEoMa8S6NT51VRpvdapzxW
Dbzf3bUZaI75LQqQ2siWH3tD8xXuBc8Tynxb3lXT6kBZhQW1S33dh+EaEi1+O3TSYJgi5peAzECQ
vD/qoVc7B+s3ypBmOw36rVDVqCFtdJs8HgNmQvHOg4RpUhgiJmM1zuvdxeKsKJG60VdXs65BaVw7
+kMobe4uen/cRHAH8GipsLzf9vk+vfSOofLKAMoWs5z72x+wxXC5GwPyUIhRUwrlfjy+6+hjx9LO
iMjp4PynaPDRD3rqtXuqDtrrfpi83PZcSISpmgdJDVmfiXq76U5xq8iZfBDPzy+eClgw2vnkqx/T
2LoC4mAoEJ/3SG1NMwRwlXYdT8Vw1zasA0E6FKLGUlZimwC9cvVIVZMTdKTOEl6LEh2W1t8bvihn
8X1yKY3nOL2FtLyU2Ek5F8dZ6WU5IhD7wEjR0pfSEHD8RGC/AxZv74YBsBEYtLuhtVAKeQJJGHYs
16252tJmjcStyUbilGj+Zzi0AKnbjiQ2sy4joaURMHRSj1f2+4pW3gdUPMzhyalvke1c5E5AXiCK
h4y7fvU4m3qcdYmoTrQU11KmR6em5RpQ1TxoGj5YpjjPfs6Vi3iqQigUUvewtlLJ2KevWSf8uURo
xdcDA5Nmz3x42Zy5qIZxCQ0kvp6eSvPRST9KKxQIbB9+HTq56Ex5dzs+1gI4HISNM43RHcqygY/3
RwiTIwZi1SNp1KrlBKAMPiv0+miz73AF8zQxfNflILV1wpwTHvnoGs5Swxo5ufuSOb3Naggx8jvQ
Lax+dsMrjl4JLz8eidq5D75wCAp59aXwvKbhdhcwB3B9JtThCZKWdGKUin/NO4xT55ZwhBO9gDgQ
VB5yGuKeJcaiGJZxPwKggOQCk80Ab8MKLoeH3k1SscGxD+KJsR1l6Qf0fVGDWgEapzvJvLN9uJJA
pt3Ap3M5tsz+imK0ASUiliLFE+QarMadzbjYEKklt6do5mLg0QcZWhZxaINsvhC95hoiO7IXX2q/
tqax+yW+yz2W63DWKpVAJshUfiqp26pTWtmlhyJV8JzfIiX2BvpNM3HNN9a2MqiESco8juGFcWBJ
2dWTYCQVZsx+fu39+4JtKxka1qH11JDHwqceA9lxPgczuDD7f1pZUVTKDHMneQDIYirAWUjowu1Q
2wc2b6DBCwMp/9WpTw3TUO0AtkZFL6WFP6G5KJSN07+ybPvdUB0aAyUVf3cVLTulDYCCsPwA5Qtq
Xcir0TvGOP4iCifXqrVqgMmBz5n7Z92Fwl/W/XDqlrAY2y+TdxI+L59t2UhL+Cg0rBOUvmkvBBrd
4+puq1o6sJYduuARm8hnZQVXSXAxVlyUdHZLmmbYR90K1Spx7qB2FyB3VnRKXw+rl8nZP540cP2y
j535ZiF8OhK1/HBVGWUVg+Vj8HP4eo0NNk80/xGbi0o6/xY9cteXqEOUviAfPJ8bZY5f8smEZk0S
jPVS7+DJjzG++kG2EI6ZcUS7hUP0+83ZKaJIKGVdOkB/JmlJm/kWwff4ZJM+lmkOwwVo3tt4wWR9
YIV7AQ6HtOX5W5Pbrj2filVU58BcyIqje5wEWLA12qFmEjf2SVTLXMdH92PijHZF4y4aenQofHSC
Gtlmwsn3CDTFeB8mxkOokK+D8eXw8GJCU5pERGF2ZYkalU9bbj3ZUBhfRElQ0/4qoejvXMZ8mR19
GKEkxRtvtmUb0M8WlwS4Ockf70nyYGAr6Rv4qUI0vVcrBRUiu7c9+g5PJ9WxKpTLdF4YLBrbUhu1
NBiuit2OUTpktACGuL/W6R/YLneBhjB5QcPMHFJtQ8x/5FC+YNmBYb4B8B8D9yURT2Qv0TYlFFG/
8QFvbfNEhQjZOYE4r4MRKnixqHFPfCHtvMDc83N/von0Hjw3MV2bdzXNHuHZ9pYm4t7efpHTt+OI
RZ+4lOcKy2z1yIOGHJBEyZOcEE2UigppVVFERDwJFOJgngd8eDpTNvpZzQpTbB82CvcnBxUtrZ0m
rWOCnHQ9xPe0ZViJjlSv8eGB8HM/OxSffCgn5DaQL4yBl+Mx1mMPBmDOkySsj25UEcpSELPcKHZC
k2G/CEGen+mnLuoyl2tZFD0T812LQJHIAT8WwFbEqzTk8V1aBp7F5D4g0iHuTG8TQX78Yiic+VQA
FfcD2izX8IMjej/SBbAipVC/cE18FoOG8cDfDeaVP90aCFQ6hpRHiAadx3NG/x6IwrQgenfx7Zl7
QSJuDEW7DUOLfPEI/+fBoQMIgPleY5X6rJuuzWIVhJW2u88IRSthSiskeRcN0GyAKaHAiHOnu6ne
7tbqEXuJb8CT0bMzxdVPOeDfPchG0sGV6eyX9r/AsvOsyRldz+Ta3jhmtLzcZG4ZyInDcRPwTMsr
v5RKb3QaqpL5jVYBOGvBpR3l6BmFV1xoLvmbDGzoKq9soQLpvBogiQBiirgTZybOr6QkLxYmdwW3
7F1g38IZax+t4hY7f1UAwBL3I+op+kfiq7qEIHZ/7j3dcDO0bgJ4o8/PPRSYfHrZTHuX1R2Zb0iC
oB2r7A0ION2w23/aXKkfmLjJB8Em1XdssN5qZMk4ZhlRd1BUqOeStizaWZ+76eYwk6sJ/n+jrDmP
MItRD4NCxR5AvORw4QIAaFZH0MnSkfbjIZ8JkajO67RDaXAPNkyW33zbNGmm2Kz8AlWVDsyxgyqn
D/KtK9S1c5rV6Boh4EkSAPowvGdDM/SY9dkCeZ31g9Lsum2wljE+vjBlrMTNhluuEc1INy1RIXdb
D3PBtnart1Jlnjuj4u36IaNqMg/0lLr7zLom+IVB45WxWH2zuxsfTQzKUngHgmcNC5C06GqD93Kd
s5RuGAzIFWGP/KRG19kegsT8GknYfVDn4Cn5k3f+786P+q0XYs+r6nyrtwHTE25Id8Y4sE6rnGJA
3ZT1MnlkdzAxZXSvPIAM3ULBWDJkrSbAS4Bv9jmLXjW9ASUcCL7/wJJQs1dzNq/ti7mi41ixexMf
wvzKWUL8ah3mlcjjFmfx2Se7u1zGAXuAOZ/XEBGBFXNTrnqFlBe7QKXNbGyhJ1keCkrVdswyVf3M
N+4pm6RbFvHd8j+GiTdtqo5jwr8CIikqTEsq2D3tCmoPJZHaccrs8zcQwGRtmN7vpyydQ2JTeQ05
+IN0phEFfd4BPCpvH1ZzraGKiiXuTAbewJ3QMRimVLtA/xVmWNvJG4nYXV2Du+UOqxIMgIS25pS6
o5kvm5BxFCk0PWu9TzdTffSrYS1gDRicDE/rf8xQH/SedBUbFuDQzsd7U5MWieklfe57w7AgNtM9
N+JPYiWh66Ck6xKaKEQqh5BZZSJttl+YYOXj5B58vDwq2rXbsB822mBmm3R4hjPSKDzNs8h8auH8
Pimxjv+KY8K24HIX+6fxLwh8jMg7GXlQpUGRx9TXXG/NWp3yw80sWynsd0h+mc5hWuPcLt6wsWgl
IhCG/WfuFUS6X1i913iR4Av6IvRYYM4s48xaWjZVp37m+MLREexifmYeV07QCscmTVIM7lZQSyBV
Ou2MmEwiMwDrKatiR16y3j78+lLSMxn9GYE3c5wgO95mggGqJbZDkU6sELTiJPplpOQ1volowYVe
xGghx7p3YjI+f/cNezmUfCEXmiYhTQLtytXvVuQ51ii6/0vWZKSmnWYsYE/Gl1KIxYc538gJrE/K
fbVe4m+PM/NdfjS8RyWQblU1WL4QgLcPaatK4SPZbIAXIz1EioiMyxU/lXONk+OGycq2qs5ZR1hK
hOuBBvFkotPhSY7ww7twmUGU4EMCbc7Qq95K4eoH01lEV84HTIt7FyqhXEdpVS7mQtq7KsgNIp98
XUIwODLWjwFzAYUF3f6kf9mCc+UEmN2zClw7xJAVwf6pfQSKSX+1cTirgDdgERktP8FT322Z5idU
BL4/BQ/29wID0Wyzf88NW1bOpQxSKf3xA52DpWhnNNVFy30L0vTnsXV+Tc2qVrTp6T3U+OlSQ4hp
M7DYhR6q5c1pLzTeu+Yvut+r4a2Cxrfb8eYomZOkt4TBKLnU/jL/fTCY9O9th6oT/ao3d0plxHMq
aJFcWKVX613yv7J+IiS4vfDpNeqp+Anguqn4iTvaOYFY15YZgDz4tUv+Br0kpbnIiV4raOQbPtCs
LpE+NN+ULIMK+8/MwG39Xo7fZ8gzFvHB5moYaDD3f7/Hz1CCJZsTqjxSWn7hNFHvUjO2XBq+BuY8
ATagaytDIOBRdg+8NiXouF315GGB3gH4X2vGyhg34M6na5evPrW2W1C4Tz9jrQBVk+FkxZ2PxPSF
h7bycRnI4jt2NZXImQyuAH002BWV2MzILkF6PZkiF8wgFLu2CtCLqaHiZgjdCHefn7//7LhA7T9C
cm0eLdDI7Md1jlOUSJ/Bf3ESmnjT7g6G54KTefapqRJEQoua8lOLfRP/PRkXzxifykVxTKWqYm7m
8gwbD8qDZcEnDawLVWUwbSWYiycGhW85PHLaCuSIuSNgMcPoGD5JnyjuXSeayIkc1AXliMY95VgG
h7Kcc2L+BJMVW1OK1+Jc3XgUFZXKz9tFzC4yHULO9k3yVp74PqjLdfOe6QK3EC/GpyqTIpNidaSL
Ywxs34IUaciEz9No9tO/dP2D163G8meoZOh1O7XbInpUpQW2Xdsg4NOT69AQeJKRlJsEPAmP+NeO
8a0sulWyYkWzp0pAdtKTLLjz7KcJkiVuLwqsz1EV854Nc1yXKQjIAodpzc7nSzwE3D0bL99+xBTX
upqEvF9956Wy3OQqNMhaqs9P5ZvERCPDU55SkkdCye75NzEXZtvhF9pQrDFZQA7sy4LJdZvSNkGm
eexWChpxMkcnnbSESMLzr+vgTZ66Ta+KQ6JQwujEujV/6r2Z4DR/2tepCa9sZVoMzwMI7U8a9BWe
74MXVCFGeLsXcIvhPZPAyjwjGm8shQ6qYEkrlhcuWvXfADRvWHiu3q9UgsyRevmuHJla4Cs5xrbN
7LdN2AEshTKUnG6d8cnRV21Tz6OPzXOcZNJ+TDpgP2K7x11LTZfHzoDUDhDoa5/yiHvEE/kQYNu6
YJmeRWi8lGunY8kAziKx1Mej0hKIV1+oiXHzfugSiZeKnIQ8Hzr9JqutQgB1HUSuxtsrJEVZgtbp
NOVRcCSSSsxXilIlv+gY911D0iyO9sK1/2kaMGjMJu8GsjFTGehPVg3mfK/ZXLTO43Jj2xeC2wtO
669Dgz6hwPSizecgyseoA7M3xClhrhEtTFgNTPK97uHHcDCjzVhG+riLyo22/B6pllB7qoeRSHoN
mQfKiWCJQTpDCmsvyN08SGfnPevt9gIG9X8wmOwCgg9rl7znYWIYARuAL0i+He82WglAncyzQm2R
BPucj4AI9BZqZT+bJqPlo4nWoRH/Ag9E8iqBHgI/340P/hN8lqPx5VlzZ9572QVY0EEmmyDXowlZ
oHgNxmWUirJaRSRw64TCqI49+p7/R9REaKBXEtGh7vmYsziujGDM2O3Jx95x83X7r4D6tZhJQ1vG
U+VG1ntyB9fbOriCtL24N8ZQM6X1dCL2k3D4FietSpcZl3iC9xmXDt7kH6AgE0sOlxEIFpgkFO8R
KK+iC0YslmC7hod6p0CBFC3BCah571XN8Yg22izk2DsaXBrHCG4Qk+ZPK3t4YgM0Qm3OpfC5+OSI
lAHfmKFwXVQYFZhISFt6ol6OMtAlZzmvXe7oEuikzfjIbe4p9ra41wwXTK82px7xPqViQBTQYR6i
Vad/OghmQmK7O9UJueCVi4PUsB88YmjBjafTazb/M0NRrDHp/JvZkJWCQFztvKgZ0eHuvWUjYqQG
FqsCTODozCBiLKXdEmCIihnY2R1Pr9cGjhWuvfw3qHDkxGW9LSih8hYWPSJ18tK/nIaweIDKv+6i
S/f0FECkljmWedluKO0y6A9gmBlqdu0noP2I1VYiIlpmiur7kaUeYtq4GO8E8J6wn1bAtm6+Bats
rH4ro/XdJCNE2TFVtK2U0CtuXizw7xZEhlkcViX1kj6IeMze7oyJ7ApBD1/XzkbMFn8U0bEM5Evj
s+RCya+SA0MtyUkdIArDX5q1JLdTKsK5lVRV1tv59uAEZFdlUTwjtV0xtONFxKTNPzfaCKCXiMQI
+3TUeNv5MeWsC1+2RxWHnJDiL3kz59IeHD03nu+fXoVTNzbgzYq1aUlIHGJMC2IdKq/Xu/PUXthk
jSYWX9CY6XvvNHuw0zeGFng+mTNdR5pbsVjCTwZGR4EWSWqVdZhsikpe6C0787lAJ/j5JHEjXeyZ
1I9+EiU0ORQpeB0I8souknFz5tE+D61ixUwyfe1JZgfcUEnJNvF8SEk7Je8OCNWOtsJhY+YpPaXy
RhBj3xHJyT2Od6GyZ9fWPQus/0aNBRIdKw4uu2SRUmsafT7pBd3I/RD4N8aPDiIggUygKlMbhaTy
jvzp1Nowjp6sUWCDZ04eHd7Cb+toPjO5c38CA+yX+UGFHsymrtGysDxhZUc0dtz7ZW/wjGHYaLbu
eUXAuHQG+S65n32+IDIDGyKiUWCid4v9ygSqgTuX0S5DZJwFCfkXXcJFJXjKsxhqSHuh0ERXItXL
qSCnPILiab5SOxMgBG3huKjmGxZov9WBFVUS1slHlcTf4uCYRA0slcaodguZQNRed8hvrmhMdt0p
brdGKGGkeYH6pMb3wMysmC8/rqXck5nx+9tqBFGaByNqIO68QDMj07dcGhA9sdlS1w17R6nBziWl
kH2e1H5ZNuvhqO8zsG494RNlhlw6gkVLsvq/eSLdCoC/pcPOEMhf1ZrB9wK4iFblqvIn2C+gdQ4G
OdGaqWVGx7HhwfMRKPvU0wn+Mw714aDVwRNr+ZpTxaesVWxI/44ARtUa9JgfkgAZGt7L3YxDS33r
lJP3fWYIv5ennMPE4UvzbxLXf+ZQmjIZfFfdXo8CBIWLOju//4lwCZPVXXjtjWbn+mLsoaROgWaf
wfPZQ96LR3sbMzvRgHH6SerAQ8Gk7uPp71JgA9NheAW0NCHj858ktdk5nOZ5bwcQk4uj8yf3OydY
tOB2IvEoaf7IEnBhIDwjp/wPwJLoqyfKWbyikaogyomZ0FNMWxuwK0lnN54ZxlIFNEVNcdCX7yjz
3Yu1Sl6hxK9KWjqObKfbgjZqPmKslnpshLWUxMjVN58tT5eOOuYMGVltlIUiX18nAAdAHEsYvPuR
poTPJOkED/BaOSlLtT0klTsXbxAAMIqNCsuVzyEmGk66RjSKN4Na3Ea78LYkfR3zE7m8FFCCp4YP
D38Y65TCWPzxGHYlPJAJ1q+tpVP9ey0IcwkjAXK67qCyK5MAAMwcwdL6zy4w5hmJgce0xd3CxDqD
/BbpqZjaV9nGyxNKDqxC7Gnimp9O0N1CZs37ES9SwtEdzB6J4LPfv2w/Y+libWh9AaeCioUGMiaY
zanZ4mlePWfFE8YUeMPendI6VwcxAACnAJR2d/mDM+N57M+dS/1t6h1ZWv3qB6c7gima2uIvynC2
bqQ/0QGKcj9XoChA041k+LyJgBhotUpGRD3J/5/cdBX+q5Sh+qU8kdTXUqUERYT623TgedV48RaE
VU5phkrOMbTlcpvHG6sVGfV1g6d1ii2f4k8NyLSKOU8bAf1Tbhv58RqU9fPym2tpEPkbNIs1qu8u
W5FMXluVQExvN23BXGeFfp9Nwyu+vkKL1Fk0Mx4moSLsHLnZwrGHB2lDCOzsn4AS0P4tISWGQPuN
TejPVrK6CcQGV24KYDbGl9/Jcl3LnD6JuylLdrg1U5PMSRS8uQg1QT2imNJx9tOfuMvAKjZdOlOw
0flgBs1HUZmhIPYKyhhZPUz20O9kKDAJcQ0bO+Iz5u8DgemvtQOM6SCz/w/5sUVbWa0azLOclRiy
J7YOaRMxVnBEheZAmW+F1yeF8xwVX7zu/6/5ToFy8sOVG0czuUIv962waPTbN9cTqEJne4Zs63zo
aoJQO4C9576TQ0O6688mOvE9H71qRkBJX4pHzRDBrxvpzQeBCe9hq83HCBt72/YVXTFsnQZYR+fG
EWhl7Jmay44YI3+hLjc2yNnlAbMjxK7BenqLUc4AcvK5Vh9dAnmgbxhE5CkZiAF0k1o+6B0aizrA
1aAD39V66hIHVgw8q0x39Gf4SFOOEIJ4FNPyPljEEUqCE5V5ondYbBRqkSDrxNZUSDseUNQExPOf
QztO7J3XniHLJ8Q+NEvVEOo8yMRCpBda795EJq42icv1dzE3DN4dXsua2pXOIAJzAQ/yYh5Ap9Ib
Iu+cimVyW5ttBxQoS3qahdSD0BRiAIe9pI4MoHCKDNCvCNPNfIld2iHNblMNQTsL3qltEd8Zw+E5
17kPST06t0hc+42y4quUn1kQnBEoBSIvjV4JDUpgzbGneCmG2rECvL4DEIgJuJ3EbUFbccVpPQzG
3KtLpMvPXv4rwMH64Ehpk7JG778tezPYR7ZX4uZdcz6p2m9eKbatLKAt64q0pytDjXINjympXG2q
EWh3eoiv7t8TuNj/LUt6KXSc3l32fnz1Ca6KR7Hw+ByhdqiZVQjkV0L+9ysWzkvHU3ZmeMbw3Myl
e0TTF5hdq+LSjPWZc19Z8GNgU1HkcA0sWQaRcMwn0U6qq9oRKcOEv0zabx2nb0gzshFa3i17assH
4sOaKhBoirkFdLlF1QMRd5zKYcrzbmToaByN+v/9LBgl74kp4GBfGrK/vTegoGzhJ0DWjSCTl+Hx
/RvyhQF1wALYpQlM3bVScQZLNS/00jeBGxEuGdogNZKhFylvd5ajpt0pfgnNTaw8WABJ1iUHFKEr
BmOvK4sUBBxtq2RvULbtE8Bo8LT3mXLF3M3evs/t3s66Iev1pXdgW2nOnYfCyHmcMhgHH0f9pcf/
HXE0dAbvcl/jSOlQvjCreAV1MxJX25tgDGy3OQ9H0FGgssw8c4ze2OQVT7UOiktIqZXq8kkp/QMs
DC8v84zoz6HLUgIZZD/gNjyk4Xa0NdRL70Viwx05KPSPUqpjQR8H6Ani7qVRSuRaT4wyrU7ENwPN
AUHJoGrv353UwoNvdcNDqontN6w/bkBKpA09tJz/Xvp5c+/nLMgpeb7yCT+Q6WQdOxwdTLREjcKM
OGv8YFi0fDbfkIhZ5kTpOTVx9US0yyOpuRfPZCP5PhTjebyRBaUzFGAp+6cfi2cAbmLLV2nqgq6S
mVzvZTAnxWNPm9mmxR4SzwEL87V5bUrvjrPODwQJDxdIeYy2o0f0r6U5SV1bHpduMinjFq7GeVFd
YVTmZBLkYmsxirKlheQFUR3nRqLY0S69V+sHhyuO1BDhGRhvWfy792opDfwbDrggvhgtcV3uBUe5
1ZeCki68sNJlpKcSUexaqcZjGHaH3aBjsHkaMiHslrOHK7QHqNwgSm9ObUUcnNSpw9YrKVrSuuqK
9UEKO8SMZpIpvM4EPsJIVfnqg6MVLdPiIELCPjSqxLE+lNVta6JviQdEV+e8mtxkr7HWh2BR7ITS
oA9eesGdwaPZGynEDwVJYYT8yD5MPkl2euAymCW41aPfMWobjAu/AB0Ow3BxaLGO/ckzGd+1i8N9
xdmhAzU0bJXcGpIE1l5OmH6sDVaMWv3bYuJEKOdbzDqTrHQPkAMpDnDfDKitQFJoS9q32DXnONaY
+1VJ/wCtFn1nPUpDVqJIZ0UxKikv7Qw4+KUS1wvT0+pxJfgKvywRlWxPZH4Tdh3JDupUI5FfTQTu
r32bxl+FAFZ+8MpcnD2csK6/Zo4pOqHHT6lVUSgCD3qjEeITPCuVVUxpGNmkm7WisBaE1cQR6wzk
AE+C6Qu6odPskLGyvLfRoyN2KP16TXUxbBT1r0dfFbC7fhnzEakKCuMCdnzEx/pRcO/fGxBz8Io5
qFtQNi30jVS3+emN46LNYabrmT9wzYftxzS/0J9H/EITfynkS+frRs5Sq4YydcP3vBj2mGHuzO+E
PhDwkmOnmyKfqpzx7Fj8I9Ixk4o9NfcoMQv448QfVR3ivcZj0K+COeLAKXrjTkJzlC51zhhvCqtD
SIMeQqUqdhBFuXOkIo5fy2Ggf+zkrDYw04bT55OMK3dOLhDC6H4xg9Ai4m0TI+NvFKSghW12c27B
bRk3TYlt8DAXlQ52kXkKdIeGddZxnM2/jzRURrIApvCG3SqxXHo55wjONgX0dNzxuVe5/u/5fldL
lRVI57OlPk0DSynMw1Xl4+g+N5840CSd74tTJnawm3EWCipDvQZIeDuzsivy9iGx++cQdPIjal4w
xiSM8zMqsxIpNJDw6dTKIDiljN1Cssxo+fYwM+5mnJqPTwlAC1E6T7aRIAd9Wn/oyC1cYCMDyrYr
OhhWuhQj6btjeLM1b8GJMrUvCs+Uk3J72tLs2j1Ekl4c+E3wVY90ZC7vzD8T7bc4Ar2cutCn3bCx
2deejbYoXqAYiNfbhU9+QsYoR8/USjTtcxY1cQ1/l8WtCObOFMNC2+hr2WvfqySRsh/6fJX9W6EN
XzxReIhqqfHxNijlpyKYzpoOMFtRT9THMwG0Fd+8qSb2meQiBbnLqy2fXfIzedbDJ0NBoN6UkJa+
hjDzwoPSfshX2Bdu1+L2HaHj56jtxW7eg2ya5yOfVYASnw+PXUHE8+dOZ/lPHDbryzkAMVRx/piR
P3FUCZqL2Z0AgxU366Uxo812UqzXqEUhuK3d9CeLx9H+yOEaZumRLPbL1XHHWn+EXtgX6M2kFJfU
7Z9diOMLDMTYFkun1L05APYHGfXuXnZPv97AVLhFoqIdilRPtG2lypLaFfnhAQeq/N9+WRMj/DTX
ULEOCzBBBnarKS3ASGi9BfQn1erHZsdNdskqFh47G07MkqMnyYqaLTqZHDn2rLuWTcQaNKGKn4v5
wY6mFvqzkI2rOuFDnj1hikeOfuzArl5FMAeYmBfgCKUUqVUZMxuS+OBpgHb5xTYhVKWKayymB2/r
XNFb9aj3ufPDqbWbxYZUiW+EquhMGTAWeC8P9BJn87C67Zbh56eZlKrXIt39n1eu5k0o37YqDJwc
KemuLNYENhQOMfvMBzuqnKBSLf0Qo+Ci6q5JqsG0infbapVeeW9Y6jS5q+PpPhd0FekLO78aJrFh
dmWrgZlVSteuc0rrcDim0mcaWw9o6bGNNQBohi3nD7NmN2ZRCfrvckyBMN/OWXSAiXGiZCUTeXGe
zN8U4p9pzkPyYBCkm6+/CsV3BmqY5cx6fskncmrnPh2XIUNZJcfCSxZWcYfg3Joa6ZvdOXYS34So
UKeGinnyqdZppUjORfcumZcbSrw7DnyRjOBqU1s9i1eJMrS6Jg87mriWxxZsKpXiRW2xNTYxy4nA
4nV8kzW2CcHgOHC1mi+Ufu9cQ4uk9npmCJMuqezQiQPDNWN9XNfBzMBYvZ4T8oJB6LnIPTt+RTyH
7asKyOmRwj7MgQRJfRglTobifr/02k8u9rhGY9IsAHCimG1JmCebgBAJiHBPEKo8qEANTaI2DW2c
pgVTM0yy46Cmbh4mCo2F4vuBFJhao5MMoJ+Z2yjLfoMCh8qRKMGxXUVHvQ8rzm4eo1KyHGFV4BO+
e9H4l4D2u+mApZd3KxUp9NCUyUMwxd8pkfm6Wd9YfPzLBOmvKetoF6dm8E6XpHFF3EEvKC33aSlq
uENScpidErfdnZ5KFVLRUoH3EcQ6dVuCkzARXpT9kL79hxfH1wog9BrDTNggprqTtLVzaX7cyL10
FsC/vkxMDBRxh25A32AJOP/jjlS1ix65TTFxVb4Psq0Dvb/s2jCE8Uno5hduou4MLMhFnx9PGHfO
cUK9kiInLnJh9aEnKNfhVH+eGLfoJrcLz/M7EIJXrAK1M680/7+kePihQ4/4+NKwxVgdZ4f9a7AI
jFs1czkgHcUqLQtQj6R+Y0nFItPZqJDHtpuH4VwJ+APyRNaZu8JyWgQcoN7iMH9xHb9nMC19XikC
SmtA+/TjYQ5aBbFHRmx/1b2UqMnR5l2HPxG1q1WeDc15kzwYQYnJIyu3FhLGey4h5/aN5WnD76yV
A+YpnM4mgwffmLvYINLgzT2vipPDu6u0aFMzNLnPk6QwGMYKElTamREiq0q16o34bZ6ODHMoEkAQ
PFTsdekFi3NAkb7MALu87wEGkuSpud2/w+HpyER9pgJMZDEQiV73gcB902JHa8jDsQgvdP2lYePn
iZIS6bnqZPZLkbdzDeaT13/1tQJmy8Xms6VEajqFBM/IG7lg7tfATsHN1fyE13fSfUFMlKyFXkxj
31qPHtxZtZo/QUatVPGWyuofnNoPoKxdFnt8rSfLf37la6c3mp9B7bQfDbsbB3nWyjjW7p/CB3/E
xrLDN+kTT4VzOwkXdrUR8vOJo/ixUAiAbGVOgT6GxZklmFWF2LtmEKVXGaw3e1e3dopCuYsXNjBy
VNtdN6pCQPOPYM8DUGFyRbn6PauLsRSCoVG8jfzir/BCpHMbwx0SdUnDwg0Z7rs0eRUkoG9tXR3K
oOrQnH/RVjFynmpfU6C5GyK/zeL1LEZ601XajW41JY7qVdkPe+N9QTKLJbXrpTppVP9BA/K+njom
DXed1HeQp3aul5M3Ft5G50V2zeVfsj4GhUY2JtrxaCiayr3CIASDaAoIUwWDCt9aBZilHiAjxdyo
4rOHE/zxvtY6+bIJstDqFGUuVf0WyTypqi8mrIJCyWQ/whB03cZBtYc5qvLB1qRCzcmG5lkZUTRm
yVQ64nYanzE/WJ0+eDo5hvmUS3F76YyE7b2mIm+B3NOQPh0HhLgD8rK3ALcePx2fxAmoES5KVOlk
1Ixmfdfk9/k849Y8YjjXdaxoWtRbQDNVdfzF+42eHO0rHFs/dhYSUOkHfy4KdqM9Iba5F9hiK/pF
kfBDtsB+9lU3FRCZ5IW/UTjZ11ONJJ26XUgc8TEyS7whQdcOrAIz5AaQjRCQD5J6nvtnH+FcU6ln
eUQxgMsQdNQyqNgvcBw4vuza3eo3ZVebCbIZ/2ET9P9FT4javpU+n/VM+YYxhv0kK0HrF4ML0dL8
nkhfSOVlYZJgZ9VrnfxPdP8+jCWee5xs2VVcX/rQ2qN1f3/zFywP9myD5ABh64UbBPC3uMuQ8u32
oMvW5MZgOuf4srwJmCNTcyjuMCjH3M1MTXJwXnQq0DEoeSdp4TV0/tN5DTDbS+22RgESAN5A4Bqw
K8OdIbpbtthME2QCOMNpL7UGduYL3DUVt51MsPBz+PaRoeL4zki28ZuQnO7LX2kNdvdas9xak0jX
cSS7Gt0AkmAo0CLPIzF1TjSndmX7VS6oumn9DBcJVeJbUu4xWqnnbbXcpHLqBqUBKpmTwGPVcdRZ
CjldnlnnkoR2XonQVDnffxpQNpMoj8YcsaIAnSSKJk/KjvNhTX4GxgKweRCx7bsfdrGtMipvID71
g7s2610gxz+trH7CGIG4T4oF2KTMsRJoM4b2S2FIvxz2ZofuP/WnjkQWiFpElGs5h8rxFJhvCgnx
Y4hdxq6Uir6XIhDlmpvbSEZdhm0VpB6s0IOOTfyEoTSArXGqNNFfOGhjF80fuqKkbz2EEPvPIPpu
HXwcPybJKf5LsLSpQPG3+mz3C2YULlqqQCBTLuMhv4ZdME9n87CvUMPIXja0BFB16oaSHrnYuuuV
IJ2FNHI47Mmo8F16i06B7LybgWlxi6IPEFDa94M7ImnNKDCTyYDDSJAE2HyekM59mVSkm0HWvYpO
Q5n7Ulr4Wtt8UgqDGdehZxoe39+JfWswrHA6CvTQtcbkXoFjkcvIPoYDrEEQvprKa2y+o4SODQKm
sKza6g8Q9nAExp1oJOuoi7iD17cvOY8GgorG2JXVxYVChJWv12bsKEgdjp6Hj+LOflh08oyhGc1G
ExcSHKKHC0wnCT5spwpZViH2duCnZ5+9Foj99jujUvJSOJm2tgKfIUH8S/65iY+i7CQZVy3kAoLa
ggl0rFazsFjeb5L94Ipbqk8ybiTArOSHytYRPF7LV0aXoS2jwyq7kEInm39kYoOj6yIC9bDHKso+
Q/sTSa0KTnpC8O8i9BTDAQTfQ5kOdpsxfOKkhm8jXW2O7oTsf/2tvvus126aFQSB3gbdImvfPpED
VXYwLyXvXZ4ItmbtSitQdVQdO425pGqlJoLBFBbd5MhIEPQRokJY1wxb/B4I9RC3IP4IIRfxagZn
n+EYGxpS4IQ9c/iKsOjuHEiD+XO9my9xHV833iGJgqOAcEnzU0ikBCtBHJAVJlBHe9cPIIeaCUte
UNTtTPm+Y9CXkrc2lIYm9BX1x5Ysg0QRkf20na2dxJNp5WhBT5G46+MNt8enMkdGhaMv/a4y+XZs
rWL5MTugzsCJ0mp6fQ6OdclY8Zy7Bk4V/lrPNESQzIhEa7J1hX4K1di28M09nDr/06yISKLa2sr/
XJb0rR5liYdiBND4VcZ+r+WloRq3R0/mw2j7qTIZL3OBKb6KJCI9W1zqFb6G+flLPLTBcOXBOwuO
T8DOXpzHVR/U/0w0o/rt2BlYyeEv1y4r8f3+Vmxns0H4ijBNJpsgtTsGka9Xy1v4GdA92YbnHG6s
OpK7XPI8L8ZLdr1OFTy3zDvEeWgaOWzLDbqZoA4cOXadiH1jZF2XcaF5HKbqxciqj5Nmd2EF38v/
L0BpfcY0u1u+thWYTPLnZjXkKDrWSPG3lh6nK1UlNUMkm56PFOQaaeSAOj/5GQzN7QmQaiCu99SN
ct9zNA81t2XvsfyvQMiNQ3r5h9SDgLHrbkfnrVa4zNK6hCKU7BrFRnpOK/MTnPlhJDlhjsCPp2C3
Q+qTCfD0bXB7YLqikVuSg8M3yAbP80iXWrmB03UznBnORT9wIG7REJ3KALmGTp5JWRazi/tXPypz
St29AccNLPyHwrI1/6ECp9+QrvABGBnIsWGjw6kcZwAbS7JNRIrZRgi3lN5axBckUyDdQz6+KtY2
88VPE+Uz/EmiV9hQX8iaF6JJQkhzHr6jzyv9WNJb+oI7b/jFczeM7xZlrnD98xqF9c2+dROaBV2B
qfodNtJeYzpGKVZlKHJ0mBrewFLP4chOgO4H5VrbDh1MGrTn5l9Z4h0iKMnC8TidUL48UV4xZmqr
kUWrbWqc9ms5IJOf+8iWWMG9ys4Qtc0z5izdg7oTpkA0AzaeZsZCFXAg88PmdZBScoIDggfylHUE
CvE1e3HY1vSIL4S6vqAHEGqRxKM1JSJ66N6n4ewcWV30EXs+Wbi2C/Z5FoUYQ486d2+7VFqiQLMj
P9HbboEbsL6Lh5AzDKhjVnQjWPPB96Ai5uskRGE6FG65Kk4dWtqmOepQXSIahchgpVmv9iw8I7Lq
jbL2ZGuHeNza2MqTVUmjAuWMj+FSSZGeHaw5gFPbkylwzJuJIJDUo39aj0rGOXnv+W81FpsQfQVu
K9VFXIJAgj5+7AG1y0KYXV9lVwuXDJt5KXxBkCT/FCRxwMDG8VdxBtNVVOrfAEQKuwqEUly9pT9i
4skAyUWwVfOotVtNXo46nC6Da2RxViilSJ3S89Mefi5Zd3ZBIZPZ5GfzmfOCBa+5J1EIXXkMDOFN
FoVmM+4mjgq0wVACQW8nuDp8Wzhn0v9E4Wdx9FkjgjB5vsRrmxnpal25q96WaAEVD+iGw7tuhnCj
fTm1b8Q7ky2E/zmD5w86wTOf7IKRbe5+BrCQChLd9EhBVnNHnEjLC8b9q62ynd6KlRyGd6p29Csp
QTzJ81KaO75WrQ8ts73euxoSAfL4xMVQCEXDpan+5TmJJSOwHp9yqkgNQJ/SpGBnnhxEHPiXSxL1
K9aQkcjwx9n2YAPhGojdLwRX7qksbRdbbPvTt6IERvRc3ojq9KEZ1ACo5B7UgTJ37cjU11dO4JVE
dnOgD5QODow3FkNCLv8kcFdK1IYJByoUYwylgNd/a5RwDEcw6TNzUSp8G40S91fOLISlCXXdfR5L
LNPdMaJZT7E12euI86BoHHBMdkCGKq8Ez/Jj3UuDBfmqClcVIwJ0h/2Qhhfz/NpMIwRi1NHeXQ3Z
/XAFBeA0eh8A2hFzcaaHjy1VR7DJGm7Qn3hM2FNc9dZa1m+lqaOQv7W+siYLiD5jUK/RAn1YZ2km
dZ8mWRdXH0f8ZcOKpj0ELAeX81P5E5w0r6Hd0iovAH+2embA6MFv2/YbN/ldkus0jnGjQw72x2oH
cCDPw3CHGjZT2C/WZJY5zqr9Bwqnkl5V0kpTmM8XcaVuM2Ydx8585CEm6hnVw0NxxLqr/kRd0/jr
5kd3K9Mdok2q+sEhRO9QWpLjbDOnRlGZpdbKXUXFbUU7KMzL/pfn6cCPgm5LwrCrRev2QgQiPanQ
cw5yEO/KSW+OsLzZIMJaFl9LBcSyYuaGHQNGvBJZJYtq2qKSxENwP1cokY5iF28z6leJIEBeYUaA
Uqn4XQiiq/Z3abig93HxWEQjNiE3NxrcbWT3zr3SvuIcRosFCVA81kUe1HP6wAbXEpPbBCRHZQN0
jdbRaV8GeFxUkTZOl0eMGKcirNKOKVWU6O1jEfleKQj6WZAVF4H0RHL5/58MqG75dDVHCCxBrSvQ
L7iep+X3nuTnAbG7JtP/SHylIdQROmcua1LjHaGEGGSJZqdScdYJ+aUjvA+ygcCuNsJNeUuVlp5w
wOcc4P/4aymNau9Z/THOxZrcDtdx6GgAmiE5kLAOgfgrXdRcp3utWvpm1ou0Fjad7eHq2eCJXEwS
wW8ox5eottjLPMRXKak/cbwuBVsMviyyFSZkqGIQQ+VOqJJGfz85ctmkmKMeXpT0beNLhNAQPP53
EBP3zu5apNEXctqzTs2EeclrTqKmFDe4+Ca/daZ9q/5M2nhR5i8HPcnAytyqk+9OWnb3B2gBLUKV
HHtrdXMab21VTH48muos7LLNm+08DVaqMr9aMCyjprsJYJVROLWX9AmYHsh4qVmHfvW/d4GC/qzy
MfYlQqKG94NDNptwUoUW8NRip42RYI9PHdlFXjhf66E0Ia3tlOPdROsnynee6s3tUTd/g/bfYXTy
FzcxS48KeVj/s+uU/HNQ/LDoLI3U8+MDcg7ns/OD/jUJ8xQ2sUs9Ipv6TkOMRM5MmZBjSjVxu0ou
OQ4AYQLZXvcuDQhZxzwLxA/OU4ZlVNttjmVUEW+4Lke1ltsL99nJiJzP+RZgTeahDrBZlrZ7Vk5z
8/2s7uoapT3ewAsZzSZlUzEutofqxAOfDwauiTGfa2ZUtAyjDvlhd0vQftrcUfsRK1wLtwlotzYV
AV2Mq3oQ+tqxsJ3kmwo8t5/svJrbDu2YrSDMew4XJPIuSAcn/cZB9FC5j6JVVH5EwOzza5tZk4bI
PKFX0qa2YW5nmrl4SnXXCeNjhor7Ah4EUmsKCm4lFl1AHmaSacLDdTF6Q/qDMWhiQktDU734VrJX
ikBYoaW4RzWSYJp4fXetaLOb6Mk5Hez93HiHoMu7AnFthPzJQzz2kjKesFNsAnHCL6xQ5HZJ5iL1
iebWdqMBkCSkHQ66DCdgal6OF20LyjnQEYM1X+BBizYzqxQ7TEZZaS0uOnrlJFvyvtmssdqxzKFR
YAUR5drKf4pqBtOBqYYfwHaEzbQrMZ6WMSKZTQfqzX+P+i4gYkRisKTffK3w43RRKVKKl8VxXx6D
fJxGP1ysrJJ3bZ5HTfN6tyITqDIF9Gj4y9i34E0cDTBPvXrrRjDqBmda/TrRztkgyT4OEUFa6Lo+
vADp3CgvM18iRRONwuVmys0xTIrklKYyUkck2XFisWYxS+h/BSEy3PFXWxIeb7O3TiGleWe/G8SX
aIncVoobpA5JDoLz/DsCSvnLzVtu6Px3pXJdCY8zfEU5aLcnEe8gGrulizrL4iXk7qoKRuJCaQcP
xCmmjB3wdZIC4USIZA2MwysqOeB6LwXPeF2577FZRpA6jOl1xZesJJFvcVpnsoNpBdWb2FDmR2sp
VvRkPvOF2k+D9J6gDZQM6reV4IuEgKzimW5/I6fXUl8qEz/JcpaY9ixL9k9FKBo2spHbfpREuIoy
BKku1fiJa0Dl590I3SafqEfDTcdFNJFGBHTJi5vLRROFpOByRuqm+I36ehVeVDuASeck6E5rs0CK
Kdoua4Jf2/6orktiICd995B/tEF2zXPpee8PWbr5Y8iM4swJUn7qqJc04HMu9TgiqrN8FscXidv4
ry4j6cMAb5UV9XMZkvf567OAT38oqTa95COIbNw6MRPVJsF3M2o4XngpGiXO0WczKtkbACqtpTzT
ctuDpsEaMtJHB6pJYHnV6IyyyJ0yX24Jrxnqxa0ovwaMmyfcbQMMgBtKUEah3gWtrduOLVwCdDeC
B2ffBINOAT9KM8egFx1V5UglKYdyH7PgUTx3OLqxXGVfskmrUAnGoxIX3QzQYx9lZ3dqRnE0cPBx
7ysTmZzYpab5R1o72zXJN/RZWdVujd8Zn8UTovc/lyRU/dtze4Y8bfhbs27ND7Xm4guz4Kx1RIEz
xw8WsGnAa/rNUZo/a7i/W9n5qSGsyflDMHF91MWWLlBgX2i7aUSKhXGJlRvu5AC588GkMa4RE/cx
ikKNmHrHA/AuQIk/KJ38XGuPw3ZdE9Mny4HSAOmTS7X7xw5slt0lvz4WaNjmQYxH6OvzoMa++YBP
EOtIk3ezDyM+2yALLji6obOarVxL/Kn8MmYA92gzGo7bXUyYgMfkS6urujHRnmNq8HyRtmZ2mqgT
uUYR1ZVIXMYL4eI2SnarB3eWwY5yIVcGLrUnzOPy4+5MCW9VLej8NPs9X7cIftOJhbDnPThr9307
w/+e4V+pHVR4QsOsCrtjE5R2qZaTfMC71IT8+c7HcU0/2vjVGDWW9uwxMOTaSQUCauvie4tzW4yF
JLy+OWvrzkgDIO1kHHapPdKSESHsHRGVsfObfwOvr9Kd3dfLebG02gnJdCqXgEFPSWbl/Jdzd0uF
s10Mxxu06NtmwtKiDwbJXZOYEKfTylTm7lOH8T3OJfXvIxWoLdjmR4Vab2uI2ND+E+vwzEkjUDgl
3o2lL/80eD/egmGrIjexXw6OZgsmQc15i2IXhGdlRuPxtxVTxD8aUsjTdCI7bYU86NrreBxT336m
5rZ76y/l/hqjDHMzePnhvcnPFDA7+tudQV8V+vLXl+Ffd2QOMSkilszIL1hcOuqw1MW8kkT8ddOb
RpUEGN0J5hvfZ7RbLZLiQib9gVUc5ZGwIjLS3coj8Rqc0y+HhQzOg/ld2nM8hEbv9lEkRxsKqWRx
7MGIehyVsiR29ySUyRvtEcLeaEJ/Cc5VjohFwgL2CevaEWUlb5N6f+9Ujt6LbsYTvtI47lmGAi8J
y2OW+MhTrDmy3aoQMQmm1z3FUdoPZ/jSRzmf4BhJfD0V+pMCOAhJzq9u+m5Rd+g7vjZqPUfbOTYs
Iutw/HvyBPFfi3anf58O7114FmaQeKQ4c9FBTElM16S0UDIKmu5ZwdXyNK9SpIaepNgiBd0dlixf
sbeca58/R47DFRiJ5apxfC5eHsGK5LIoddy76WQYGhcnjInduM8qlRHDPJEHiU3SUTTMbKczzzc1
4/BTs5H1aFIB5HMsMVithVpMm4xBZrb6bZHPYYcnhMHgAg4aq4nGybaVgIHxl/f8YfYfuzkYQMa8
abv69y8FcjmSprAqD8cP68Uhv+MO/4zdeeVmi8sYhcknSxmnsLVrz09s+2pWOjhyPtgVEYOyBM7u
pNVvhIkYlTLt36hBcFa7viQKZWwBXQ5eOBVTWDpmGHJvCNJaV6ieCD+xjvazKpUZ3tDgP18Hr+F6
GWdTJqhl2PBQYd8H19JWLFXrcSLvb72NY92weMKt8sF4Vj7ByTxBE4Uw8vcBgzGC0AXwVG7GRyiC
zqvuGkGS50HVNn0u5kSKzg4OxfdCHab1lZD2iDPoOAqurU6eksZ4oQn9fIeQoJAcUqwUzRWcL5LY
NwfMwwR2tU/PIz9qERoiNapHOrEmFf4mDK4x3iEMlvOOR6w/3l29zHAfA8xgN2AJNbjOUN/MbYaF
nFY0AKAKi+8MnIobajHAu35LbhLGJY4AT4vmN5EDlvqsM+oG4OUHPRt4kdxAWa/scHffpfrGdzeC
gOBV5vfrlJgCWPl1JOJ7LS+vU1wmpogxGb/uOJcYwg7PaELDtSytejwc/NXtU2A56jm6GGnD7OLt
WtUieux/d8vRxO871zr2y5kslLZHKEROdBNyzG/PsCZzxNnp64XaA7QM6cEvLvh+D9VuwVPezygD
pHR8tXbGZG8OpLiH3CbTg9WGA6ZSs5tQQ5GFWd2/KOBP0ymQTkt7sn5p/F4+/Bmg4jl3OcSdKdK/
3EsldJ8kcMFC1nbhDwkHEUki8e1rjA+cC3elNZSP4NBZcxX7FrK71WBlNM7DyoJwkuDS3qVsiDI4
2bIzit4quja464IMLnOo1wwcZlTg7xT7UXRAYCTkiATthgX/TsGmgL5F+9ZWKgejvFkr8L6cbVi3
j49ufDeGBNdgXlt73aMyMdHMNd5kSbPlf0D6Fkh9Thjc9FM98nSVS5+l7abUBKWKP+0ZOCzHuT6j
LEwlQ6yMDybgWNsw8ocqoqlgPh4HG53Y5Fb4wNN6pFXRU01zvt+UJGP7dfvV1xbwfWaVEK6OOfU6
mrq2qYq47e33ZwWympknhWVEuQ8blFKlnHSJCxGMtYAr+w58IuCkOp9gVP3QHz4vLaR3Ez/LCzTI
/RtkehrEmfwOX6AhOMA6d/NrRdf2bNEquHQNNM2Rdi1FMZzB8sKlXvLnIm0z7k2fFPxGDv+GdWAa
LoUPTP2xMMjnZ1TKXhTfTPzvSSmCZKuW4rkcElU+I5sXwh7mIY5oUnRLglZSBI5xlTgKstStD5+B
v9a3zzX9o26GydSDnRfZS7Jr8BR4unfV/pwjfNhX1AjL3AfLIqjC3rCHLOeqQ5X02Oe7PdTuAhPP
w/V3PkvwFXOt/ZBHobEw1tolhqptjNQr5dPGHVMDFrD4T3XT9a9n2eFbdUBg3AdZylPfiTSp+kRA
1oAZSKCvH+PscAcER3Lnj2eyX4nBSG9QShHnjBioC0TQGwwu7HlkFYNszxQYQKA7LOUOoC/jiaFn
8TZCA+DW1AcUMT4KKHQG3J4ZrEXfAPgoLftH8oX9CqOy2HPG7shyMUelpPA0JJJ5b4Tb+glW+VtU
5854QNa3k3dTwj7MwP9MuMRyj1ktPPVioDeFEQGGDk4G9JIx4zxDcg3s8NcdVueEm/CyAiaDODi/
E50yP+HU2IIzuJCeMcIzgzPfN8Zv9U4mK73InGdS8pk7iKBe0s1NdHZy8W+z3LZ8eUMueeu1+nX+
p4vus5Jk5Imd1UcmqR72PqTiK+7CXbu3UBGjRQ3EIDg13YyaevShj5otE7bS6wqIsW1kQp0rRUdF
7b9PPWAVjR4iKInxxkQO+A5KWcwQIPK/+pNkiTO4RRh24/WkmdUcAajWKGZO2RlAl8bKyT8i0VR/
p43feqjXeGdM1WgCWtfuZS4TeIocOPBdpMpMmDZdC2CB/lTiA6CbxWirowkCcvakvk1q2t02OQMF
KrWauN+gEmOXCFyvvHd2uQ7NCaF7qhkFdqdafxo+cPrugJPVXC8Qnrh/fNtL8zDh/3dt47AcbNaY
B0v7LPo/tqM+VKsPyd6N/3zvlAVfLrIe+NjgCrbpKC9NMLbcUp8nd2ckzCOUIjdkC759gtvIdZ/K
L3x79i5REqjYv11zQDj1YxAMhYlNH4L0wFA1WMIzo80+GqtOJ0OYgpPxIiUFBTDZJGXn6uu5o3wW
hdUIdTSpvWm9G2cg4jwTBSFWZk99MtmLpZ7dltFUG1VYJtt3b4SPxHbEexO2wUCYJiULQyPq6G2Q
XiF1yxkvEhO88wFo51K+6O0tNIL6+ZErwCvCrl3ND3Poci+hfmXj2jC6XntfZpyERofpeBH+dFaF
Lx6CrSpGpstlOnwmIdnFNnJOHhiuBh7XPZQSjHPyJ7O3ifaqu8sBgCugD041KYYNhdcKxs0A3w5m
wkW2/WEduQKXiJ+1lQ4oDJnp/Gqw0TEgO/JpKqkvcfoGbcghhLfQaE2WPu3X4r7SbYyd9EQH2f4S
wuAtECq69C5eM6xreCxjrbzPgssfTV2aFfeYb519R+5wD1UhhOz2nNKS8DVvkUQC5HEvJd7rxyEx
c7I8ckXVNOU7uP2bN70QKPgJIp3Er92S1I6A5R4LKufSzVZUfzw8w1s2X99UxLt72iPbZrHEEWVV
zlrqRlwaRvFuAMbNRycGKNP/9DIUf17gufZ4/dH6YxYQgB/FjnT5rRJ5llB5No+ctvZQxzrwykeA
cJeZc5UEwRAoXW9v1ad86Qv+TVPlXTjN9sCxU0xHswu9x4yIyBBgQdEZPQQ5LQDShJgi+SU7zJh0
NL3pJEqRU2+XQCyr3lYGd2bD9XYp7zscfMcobfm9lWh4aMHzcDhTud1b5gbKfs/1r+NyCFroo5EP
+NX2mUQP9VEz6cNvHj/nkxeDNoiK/3VVKII43J8LKL3fc4uB0kq0HGz6Ff1VFqfjZ83ZSc/KD0Mt
geq10QKvxhQ9Ao4wdYUglmbSa5IcamuWBWZuXVqs8XbA721QEYsRBwEiD/M1kWJENAueDXvZ5ZY6
bNK7hcNu9WlfMT1ocXM4kJ4gLqN+3Ftp/k30b22pI7+5aWAxa3os5bYivNvRxV71h4pUaKWr6Aft
DZW3E/00anHqIRy5A4O1Fy1JvBQMLVqtc3Ea53UB6y08/Xf2aSkNqLBDYbGboFWxkJtFe1A3pxGZ
SJpBMAb6Ut7k+yjqURQ0frsoW4eD8KwfOaLRslTPnGaOB00QSpFmg3Gx1hFQmq+w9yE+9Qocrxux
iloOqXX7+nCrNx1ib25oJxe/u8b7jRraDqLgD/+xJb9/L2hDN7fQ0Li/HcBw79Bnd9EwlJF787GO
FdKQBG/TqaK8DF9ZEK4jMnvRMZ//AItfj8HuwmYBKWqlMcWVLH8lUAWG8GS5W1LQToUinm0EQkgA
GDUAxFK6/hdaKS9PsaGZC7mmDZskxol3xmDc7lUYIaTOJpG6XYBh3xQy6Cn7E7XBcDcHBWy/vLcV
q7nai6zRbmJjaUPHogyp8v24cp7lkHGmmrGmIg8WaXHO0NKAZAP0u1nmnRjZ1vdpEIlWtQl1DBGF
O4/sUXRybdtGnrqEs/AFOOfM1P5xufGeGqbghcXVo2IMEAuGBTEE1sI1A3TJ3XbYdBFEPLVKPwzD
kf4eLw3/UIZxTkqcTQMlALJBXQ1ZptQRZAViBVmA750uv73xphIIO+kAVqSjxfSmnnBbv6sVzhbp
8s0xO4Rpd+zxdq2wU/GqeBO6Jp5MLF65lDP/7FHVF/7iXzqLZcWAuY3hpe1fiXo9XDbWaogjYEcN
pX45gZ+fSpOv52uF42gZMrELsEfJDHhyB5/BhXPp1iMH5KYnwJSz+ddDfmU8VhfOOm4oVB7d/PIl
epRI4p3tCTOGI4Gg4J3dFYglumHKJ3JP4WWbK3zwpFOun3VIN+KN4NQEicLV1Jws0GhgeWBeHBHq
3Yv0QhouqJ3WWe+z7hEiPbBmQ68F4Jfq9j92yS5CrhHh5hy9Q4KcbD8IKDsvxb2G8Tw+BjQyrwTz
qP+E+vIRHNPj+CK2PwHZYAqakP9eYTBdZ45hVC791JNLnYyavtf+ZoM4CeqXhs3otbyzUKScCGV5
1teZDVL5ZZtuRnLDKqXqee3aD5q07K1H9rB8qK6vtztF0J/rlRY6O7bzd3H6vWOM2KAh4isnQJsP
t9KZfho3ilwaeLJYho0i3ZPWFiEAhk4Acgt3P4keO/JRT2XQFLxe9QrY7saqbQ1f4OOMEp32BX5A
JJW8LfZOTCqVKjD5kDeHbuwMEA3fR4cLwXQoLFHGZZlglMmhTft9zzbRzntYRMqoVqy6MZGM2KS0
z4oh5WUa/yMizqTt2tPWWV9LGbJHnLWaRqHdo4FkX4A/0FCJ/0mQW0FUkEiO++f7NIK1MFQorz1J
e+tQgZ6t+mKoRCIgQAIzOKCSwedLLscvOu20ldJito6/th/ciz8/dXRo5+JxBOmaA9L01LzUfQO/
Lp6AU4rITyOJhtlsB6SvnO6auBaTpRSrBWNlf6/Oo28ownDe5iosjYiZrr9lnCbe7jKiNXpVsGdP
2KA8/uCURpIudsKCBYzxrET717iWmVwEc/fvpQjW9RO+VgmMVv8tL6VepSb+7piH1Wl5bmqdprYq
noxNuQHMH9P4qPvR7G48UGjHXnucxFjNQFlZ6eRyi7icAUGUct3AxnI+ruT1cB48gRI7N1jwGhog
B7A45/ZRbsPOBcdCogqAAwuytsfp0clieF6csFDMQ8DOFeLT0EZtDQ5z9P0/HZeyeNJH5EEuFuAO
We3A2WCpPNjwXsh5sYOqfRcpn8x+vG80QKyPfp3ivHQJFoRuVLsNKQt151rd/lDUnwAq8ngUsWlZ
RXgP9UQ3G+T42eUpXLSJoPfAzJFtmdWpsLkS9sJuovuxpTAi5GDGkW3Gq+tYtiuOO8wzfvOUxlWL
1b1rNsLgtifI4P1v5pND8q7S/WprE4zGFW8AYP/9aqPLZStetdAgITaCXV+8ta6nV4gpGOu3uEUx
gP8HIo2afGc0rNP9TlV9TlhF6OEYn3Spk0yA9b1lX/oBYl/F/o1QcA50hpP/sdAwDCrDtCZAFb8s
H34KwFGHSQbHuY9GyZGnj15VJata1YLxcqgByR+/Yhn2yaWn/XfFzg0v/xXAO7D0HN2b8FseH9Br
gk298g3xCnY7jPSovDMTEa12seo8AmAF1Fft/GBzy46f27vYztRjqkHmYC5l8j3XXNhglPD3VUTH
F2hOBrrbP51ch8L3qCSBjCWuGbVBciIU3CJ/68J+PmjsvxIy0rHiRVcdYxtThu0Br7a5s4NiyIjT
GMPCGUWiEpfpgPlNlNH+0ydlnA5EnryGHdS+D3FPMPXrJ6rjMlIqI4HW6oNfQM6QByb7omSbY3Or
JFoKhBW+XKIlndKZH2q47fHAtViXK1K1T3YD8aFLf/O8spNefv482iY4RSs6jtV/y+LDUyL5Oiz+
APzvJQyjAHtvOrXdpZBIFEJb848/7FvFFR2Vh/I5uZONStwFI4EZxF6R8yS6Q66fwZuSVC0OqAAJ
xzyVuz8bNzi/1zq7YiYZik8c9roxN74/Zd525T5u6CIMj2slWPK90uW5wxfK76R6FApRc2DBHz9J
S249yNkUsc6fWb3fIWMANcOSV1ioXjGq0vBKhJ46C71I8ArlUpAVHG683alYG3nGqFRXRJvRZQYP
PWenJxtsdP4O5g73+eTdTYILypE0M5INMB2XdYOkl3w2SG+k5A+lEce99I1m2SfMFjTvf8Vd37g8
bnRRuaKsL2I1xJVBtiu/h2H3MGml9JuWLSZq9h7IxudvUqzZilIk9K9g/iN2OzACPkj3C4g6UEbf
IZ3nIH3RQYH5vrvJ14Aqd3z/RArOxjsLpqBLKq75OC2kksy1i/IC9UERXsXK0IQacBfNnFvRrBR0
qF0DaKj/2fr18dCGi8TGS3+06Rj23A9eeGKq73mstFWQHAG8lQxgGZFvqjaxyiTJDv/bl8Z+n+8n
0vaqbdNzlXYNuLNzCRfSJSqlA5Wb0JAaa64vMQxJ+QivMeFuc6iF0b6uelXMPOczepzfq0p7H4c/
x8ktu9hlQPMLA8tQ4tEK2qrK2oG3wx8wku7vTA4Ca0ZmxNLtus26POcpkH0z4yRwaZ9vYlpA8ATE
qaf/QafDXNS3wZSbKv4312KoUSlsLRVULFPJvxNy+MAWCVU+/pKi1RhqwTv/S86vV/GT6aqUUkY+
Bia1IZUAEqAZwmVvfyJKbF84xgnS10lw3m40CNzrlPkYCbiTIKZ0pK6A1hcu5cymcasBrqixCzUT
mysrrjoXPw1AzfG2S6Kz2HpqeyQlCOUCuiPG4zqBSahv8kI2+XFmkTKHZvf2GTQMsobbx6rca0pw
dwx61D+glKmBkejbL/Um5IiDfBkoM4TZRSxiYb/WaklI9ed03rUfIbm2kjWxKv/Nj3CmkT4alz9O
NNy2imicIsyBxJTiVst5YhyJ7FPTY0y+fvlT+j+ZOxMPb3gikUe89LUfrSHK3jMsSh86uU20l2c4
kGsE50g/6YuzcyF0pNzzhTPP2H2GCRNZLEdR7Ie2MLB4SUrlU94fUIQt02lXz3A/ILiI0Bp9xn5e
18Y5ifUotZy4JKpe7ugZdQNN4Fw92D/ciZZRSc3LLLrC3LioVfG2KNum1fD/dLA3TPTgFirHFcEi
vRwC/wMGtrmBz2evelv7GPdu2IySUJYZMqOywr9S/SAF6aqiQiF3BhKrsV61lAcW0EDVSqkXgjrx
88CX6cTjgDRMSNnNosWDqx4wVD3byWfOVQa+WrNQklCqRqj1YP7lPGJW9+r8dTzq/AN22HL8Ieao
FXJcatM1O6mdPfWrOkVqrIT0upmacfC4YUlrQWA4MQD+Sv8hEzTyOa6wsHcW/CMjx6kW62AUHmB9
aSSGyVqx5LNj6ZXQc2+k+h8otfvHmoneZj3B0zxlWLi8gzJlnPakmx7Xmqm5lBVfTbE20xHAkkQ2
+veCKN/ZFzDj4qpRhf+SydA1uXMQ/OHp8CA9lFKDwHgAZCJkQlfkAsKtP3owqNmMtcB6T8KIX2df
JzwGVlxfUbboQbfCtW5u8i1U8tO7ooNZhMBmAe5KcOPfI5OlwbCH8JqScYB5DKn1xRdM8Z0UcMEF
wGl4eeAcUuCYHiP7vyba9zdnyfSn3574DFRXmxVG/RMZ5kareGPwV54RqP9JquRF7BUqrcgOYSsM
ObCPGsb/50EFK6dC1LbtJCJZQ8z/RkAZWl1mm8QGs2+nsGYlwZaYA2cCRaEVXgcVL3m4EE88u1Em
SKg2qTRfjQBQxAva6V+6Bmc+Ofugfhfi4bS3GK8q+7DIkNHbWSPV+CDnHSebBhO5OGbdaKkb/Z8Y
o5en1z6HyVoLPjdjOcrmS3GvvKJ80jBVmj5zX4Llo8PykeSLFCd5ddT/PyroYvGy70mTre3zNDcm
UUTn4eOzcGWWzuMOirewmDRMMzK4hIjUpcp43a/Tu3zAMPt8u/8AcnxFpZo/cPvCDiT1Ds8fgNTA
TyspItvi0bG02t6DStAYS5qch0r325Ghd787IJyKOXGZSyQ2VWaDWUrK2iJXYrldvHznG9iKXSP2
3YB7s3cPL5yp5/I5gyntJXA68881/hKfM6jSpR8IwkDAiF3dlm2y4HZDQVDWdwq1l2jmzM8cweqe
/rzHgNVOjnR5G75RHElsQQ/d5gmDFEX8iRWyq63jslktZcqVAcah+IWE5w8lLGUj+7NZAGrgYw3p
sEsJsOxqwP3txYvTJkj37YO7M6Ko6D5m/77WGkdqOgN4/bmYdv/wsRpWe0JF2nTFqpZfLKY0CTlq
wrIR9CNESNXAnYXtkZI0PvUppAHal/gzB7+DaZhjpd9vu487+l4ByaKFJrTYw5JXlcdrA9XC/v49
SQ03fOEwzkz8Tu6sdgkeAyVr72Lk9NgT1VmbzNmAwG7mrCYHLfIEC7HJhr8cxCckvWdKQqSesK/K
q+itGw/JRcTfs/AnTCDm27lhkQi91Oyi1BtWj56xjTptZD+kqjYsQaQ2nwPAACD/qO0L6OoM6Ulj
x2v1Xi9OUYrWJUvoVIWGBnVoeTRR7uLohs+7+ZDGPlWFdGf1N9slu6GwfHHjxXek3YlLXntA+7Eu
O1Mc8uG6cKs+2uCAYVHqwpTbvv5STqdJLrS7eoWEJUtjPwWkF/2QqIge6D6ihCb6LkeYng74nGPR
OOBjMvyMFgjO2NAre2KR1hxGjWYLe+alTPu/bTQs7M1KDQo7mzNIbISyFiy179NW6CIeNey7VWKO
w72GYHT2XPnJLd0ZpuwGuEFFIfUZt7s2+sx8sjs0WeKIweK5NLtdMercRhuTOrnpmKAE/TyztFfn
+RTuH6MswdPS1bhigJtW8EaxUJa95z4cYU1oAU+B3EpgwDhrbDFzROVAW9Z7IAU26zgaTM6Xv6gd
/K5BNdww0KIyZE5NC4lBZ8RlpZ55hRjWgAfFIEJ8YadvF+vK7LNH2lKDqc6S9P1Qnz4U+zUZW1k7
Y+VoJcQMiy4W2utmSnxMwCoVacA6i3EoEBGYmEKcwCReyBAx6Qea9AapKzRDNmfppA7hP41z7WnF
sWweAKaRAz2b/B7l1+Y+37b+s5G/2/0xpqg9cYL3Vr9OA9HJln8ukXGEYA7/gPglw28peHW4kdM0
BiARuVUIQIywWdTPYZ+2o0agjEA4e25TS8sSqfYsFw5r3iDKgslh+L9Y43TLbySeeg6qwTTdu7uy
BfsreZBvfSU7J6SO4PkYPRuiUd3/zAa73znYsid0IXPuXdpodTVqS9DTb0zQEcHZS9PzdLo/voQe
Ra/qmHyLcP52AxMYZ0bvcHBsd42KCd1/ez9eylRqlz2w0UhPeHyTlax9fOp7YlIgwa0p53ui31ed
WTeyK3Aivzqu4TyYzkf7RAFdUA6dHHbkWu2Y9Zowp4/431mWvFNTtb6cqDoKuf1nlXpIiGs/Y8iV
CWVUTuQqadb93RlVmJg2HeV1lqXeouWrZFxYZfP4GR7WAqFNCUvMe7oLMyaHld5awfAx1WL1FH55
MbXY7W+kut6Py1fWcHenwnXzpz05wqI6OUmGCcUUgm4eBjq42Q89+41OOvKdXpTyB2aNVhCbjK4w
/iE15ctzKQdXVlnUnUTlC9neoCpaYswwyZwjj+3uCLfYODyLYPVIMSBifzzrHu42obsELji1vDMR
hEtBPrsk1V9OkMiO0KMYWqn/pC6w0lFJOTpAsp3pWSvC2/85o90E1I28si71Y4LO1mbMM/XQGoge
KYjEXZlBGVS6EetyP8Wsj2tqoz2V0PYjH8xFWFQQoZeWLRTO3TwRECLis2CFyYU0dIIIxR8K89FF
0QPq5eljvPzKtGsn7ZyZDJIvBhljsQb/E9vA+5NTRCyoND34gafYUEmLpiX+4LghtItVIh9+SgTN
Xm/N3+2JqnEkn63Pro5ovS78Q0tm/YM98mXLLKFuoLOLJbtVLF1KGALNmvOHScWoCroRxZwlAokp
iTTYDvUWWEs5R8wLxwptMYJX7NuU6CS0lLlo/PPtPnOduT3WhTPNAZwyNsyXhWUJBV42H1a/9REA
5P4AEbmqCBWQhdXXe2dMMCN0Elt9yjawvCL4QkaimIxKpebEVrOFD9a/M7lJHIzA2LTod3ITU+da
ArwHBrtuPMTDcMKHub1yRbktKM89UuJHaEynKtIXzgWuv3uU/YP6tTx7rERWXwS0qSSWlEZliU+L
iOEch/hiJiZBLDE+RqA5VnnEe2kcSoGDBopxLniNL1951dkigYokFsIHki8Ex2/f9b230RYifgeD
2hrQa/Sak3mHTARgCmMoCaqPlpHQOdK2dEVbGSe4SkPryfXM8Ys6xyR0kkAftC4O5L3tp0D924tu
B6lMT3t/WZE7MY56wOJEWuB0g2BnplyakHP7p4XH8sc83d9t4ozUyLmNtb3oYeXWaxeAhYfrGGPe
MITSDancIWxGo4rGnGDkfV9ZfjXotGDLOiLjdL/HDh/3nDITFrCPROg40nlj3VVexHPlO/ViIfFR
Q1fgmqrVMFmrOCTeDnpHCHpvbLPDdd3Ohxbaf18LRi8asahHWesnFFvnO88XBNYxm2X8jLM0dvc6
sw7X4ZHDBZuXLstIv001kRkzca3gKfhHYkJuHRmPtH2iGfbgwhNk1drFKcpE2NUGL2Ix2bQICkza
5KbzwK9UzvCDILD88rzY+rblPUCv2sc007SL+OOUlf7it5pg29qD3+7uWhPJw307p7oUv0fvhINs
a9cYWLqOMAVOK9GVb/jM3FcS3tk2sEBh0uVhYmBhc69kK8PZnvYwjLbAgLje7ldTMpSGZfZdu3aT
Hm3TxM2urpm2RhxCaMfxnpufq8fMHmZ/B9KDLxbqIyv48e0ENddMDADcl/GIOvH846NWDhPW+qfz
HrSQiss/UM+LxHvnI4sbS7GCoxKrWzw6OL5wPIubwNmAqh/59v27HS2uGGhUYqkoX7LQ8zgPNmAe
x6acIeKbYUGISODeuE4U3781ir6nrsAbHNLS3Rwn5cDstYj+VvSIfGQA9/QFbnxKuFVNC2XesfGp
t37e7ZqQg039Z1dqXHEQO8zwxypLs3NNOzBsxYt7B7ZV/ndMhfnAMJvwLzkkTYCr8d3012iZcoGS
tHoJ+jw6yava7fWAZOjplByNRj/1wCDEopD4C4OJX1tgbdoen0GXJeoFMR7F8G5GogWLT6EUbyxU
wk7831t9IvmHmJs56IGlPGWvw5cwHqBd4vxV5WQxuH3GrTwMukLqpbg6RBD7rCmq5KDbdl2Zi6ly
MjIfJ6T93Yxf+wF5KxKqzZ+boiH9/SsoGi0uMXrWGKa+P+HAg8EzoamOL5/goOMc4GOVa08T6NVP
vKIhP1KAjFAI+hYKI0sraR3+/K5HF1GGa2q9XIwrtGV6730uKihNN4MYbJJXOwMofNWbvH9Bxnq8
dMPSfe+AS+vjqMOPb6oZ748Wj+Yo+iXpos1lb4acqLk4zlV7Q40fsQBPj4RpqvVymz1qwmsIZrbp
mprza3OXrFufNjZZ6WitFr3wrdXqD981z38fwwLXTR27bhnuh9+MKD5r9JhJHxndh06I0E4Uy95i
CTcxI2RQ5Tp1BEWWgQWfXfNHPMvWvkvCOxZCWFfa0zhSoGjcCNBUFEEn2L5T6+5YM797g44uV/rl
b90ddPkNkbPJHz+YlrrdLeJ0TNi2nmsHiWltrZf0La4RAnPaqi8dQ92sYyyhC/vVTjJf+6xsmlzo
J5G+JkXReVkFlRZyqCH+aylt2WcsdtrejtE5mXu2bLII/mfDVvIa9xkSpN33HtNh/Qm5Pq1Ny+fH
lp/ppMJps/tIpx29+jnniuw83F85KtBl5fTMbb8s+7Rcjab/iTeXdtmKE6vs84/WdDPnB6Hf0YUn
8axGX86sNbFwn8es/xAg262qjHqm790hJvpAFjDiTfg8pPEElOF9/GHYIdJ/hEpwt+/07Mw6UT4p
OIQc4wIPCuBhTUhQye8jR9SFGHtjm//T9j+f5RWVkMt8OLD6eU7jQ6rY/xTrLlwg9VL7/vVEyfam
uZKUPdq7uD5Jtt8vPmRzHOyjxqBEn0Geuoy6fw+MdJ91zAq0w5c44z6MaUg9MEs2pgnMerLVIqEI
59raufgz5Ld1rU32ZuSFnOhPobxEni1w0k0Ysv1YKUfnCm+iVFh2rlA7NyEAm74PQNeUeh1d1NO1
iYLrSpLgT4311g4ZO3rNfhTlWctmwm1BvaKHNTyb6pmf1SHdbKfcK+Coos/oXwhkJe3jRq6MfbCU
F7PzGciBc1Vi+FjVn+VzPmKVzxJ51CUgLtd159Qi294nV4m69TVS3Azs2wFDE2ykGEjOxIM3SdLf
H/wkzGPBRpUjJYrIln+UM1DvunLMkadMxKGT7rToUP+b84IFKcd5uvUGDFgTu8fVzIIQ6PrwFfQI
zvHmyzxlPqrgDmlokvTdW98qY0WKpgPPaPUJJmbL2o7yNtcgP82IJhjdpX6LLqiRr5AvceakzZuD
nUKIXnv4J9EcGGQt6nkZTZZ6YswRP8IuOTORXPrkBieTAQ1F20CJpsChR8FVSAnXGzWDqf9PTW7u
WTZuECqbLl6ILZx0lrvyw3RO48z0izl4efiE/qYLUgwXxn09E899fQ+um98b8if1kfCfPqRU9adM
4jFbvjNTIUpEdKv1p8npg4g6KqWQTzWhNdf9UCgb6oeW5J84Vim/cIClNc9zGgTCjM82z+w3HFgw
e2Az2ZhqsRi+UUymSnilO6Bty0/wbcCPdMqCxNyVZt61eEgunSIicKMY4wqz8MJj3/DBK+ltnK/p
7eFhT5GOXfZ58LzYwC4r9kX0WAtRKVOSnwJj2imIjatjxXhj4zpOuUpFHqeb8q27MdtgZPQKu28B
TheZCYPcrm+Lr2xGJsdMLZ1miSzAroiMPecC6Q4u9wWz+u97Ae3/hhQweOD0o3miwwtBhzAJhBok
KjM2WITVNNHluLNQ8eXAUbx1sZ4uuvoN/Of67XAMp61u6/tTNmn9rVnvKvkxU2LX03dxp7LzdJ+l
zzooq7FeFelJOAUHdeF8DDt1l7z/3cJRjgF2ltufo3XL4Lr5mvHNcHkQvzkEast+IWqmnW90DTNy
Lz0ZHLLwaSZBlAMQaU9dachhyjVrKaEXesyqcrwsJKlHVRWbKTclazQzO30eXcUi/t2dxW49AVZc
+lAKGgvTvNbApjJMvqDSGhXzDukxBoBbkcW2HYJFfA4eiNxS003K2KV+TUoN5bsFfeBstvIkqcIh
/8svmn9f98tyR4z5EqUDKdys02LaXavZbpByxrzG3RhATyut5tKOmSjHhaGYRZ3uiDEaJUdtUc4u
+1v8Gur69E2KgyNxX/mgXpAg19JcwMXSLFsTTPveEj4A2YHfGNU4+zbRuizaRABudlsMG2Njd7rb
L9kEyWZXuGriH0KDC5NE38gwztzaLvjkyRT1gIrUe/xmV/ORia9DE9/KdvHq2032QEbbZE/I04Pi
undlgA0HeVp3fI86ya14mcH9zO4kPRPL2Y+BVgWQb20APKdebI3hnU4z2aULrZZ+9KwLXieKnbRF
wGa4qhh8EMDyc5OmLQEHYH/LRQiDQVWfix9LY/+665922u//cQR5QLzq68T4mgIlYYTrdiKBE2d9
AUbZ2B+wY7RnuBiGkTkQb+hva/3zNtAYCOMyK7z1bdRN7WoOOtvJjKeI522+oTjeq8zhBxN2hx0/
3ZYO+uNxorbDVlrHJa/8xbs9Ii7WDRr5paW19qjZg8gFIE1mRZOnGvCa1e9csJE+r/2l9n16zKpC
f4pZKmyKkf3QawciJtFEG1clybYfEK50rVVKejzChJHvvlPMyjhu0fz9EAG/yqdT8XcCwJk3EngO
2jaELfFdIjSWzvcfdATNa2/gr9K/8wbt57zH4B+xVLKuA3DWharv3/p0nfoSmXVsm0Q98fxZi8Or
51Smfjc9dlXZbfJ68LxsrOfdvukPogRY4v2yUCNIO2z1jH9N2v3l7aoJWhh8vuhf5u5/nOesNN+e
Xz+l3CunwJHwYTxTFX3+9zd+Zd7SU+VgKPf4CoMxkqXzTZ/r7rdABHtDPl0woy4rS1gK2E2OWiKE
HDWkR1LwCbNSVt1zWt/3JVwNGWvrCTyLXJU3gw1OMDyakQPzEz30GefBe9nVItdbtkoiH9WeTGpO
voQGRmz9y1Pgz5oM/Ow4PuQ8gtLxYfxH0ll4vWsj2dVwRb6kT/PEtX9h/FZINWVxPZyZsmn6zsap
Dk5glcmipfh+xNNtxLG6s/hZ9mFf8f/5Ro3b2tSbENXAQJRgKXrSkqSV+8d3fdZpdU5FC7Yqgbz0
ht18i8rImRaSgLF/Y17lScWqIBzbu7Ll7sJeRLFJcOs/JYo04xj/iE2QUoARNLbO+sAtfWnGo9wU
A5OJwzHbmkZlYFzdnZFZz0W+LKUPKkCi97ACa9XzeoT5q/3yFAdHUrUnfJwFXXI9bMAC55svQnD3
utRe1Wwbo8y0BfCdwgDYcvXRxeXW52825md5vyrmrpFD6ZttKIa2HwFXPw1tGZ9urn3Vj2BJkyeo
YuBWBOQe44fmn15qI2f6/m2hHBEEFhc+AdialEtEVLzzjS4HJGfxRY3Qj7s/Dl9Ca0dJz9FYdEYw
18D5GfY0okK8/ZTpA8suPRVlmwFbAFyn8acZxwNVvcQb8v4fjNQo46haV7qHncqRyk/JWTVOK1BU
kRcGlWp284M0sQZB3Zj1RvhPbN0wZZcsDF0y8DLHnMXeW7VvNI19/8o6Q9lx066F4iO0rUvjGgIl
X8Q25XuKBAj1J4/19ITytnRm0wy5QrulftpNc/G5+mVOJz8KKtpy5ofYGXb4lcDsdR/IJj6IVIHf
2WORlZQu/maiDe599OtIuN1yOLLK4hpkO0UnSgMWDQC4+Grv7Qar04hGnwGAileG5/FFxPtExOO2
8m9uTMwk+NdsYMb96a7eIpdVdxOz6Cg56dSLZ2TIB3E9PrnGxUdnlNncUJDGWLo/aQAyMz8ETxwK
HQUxhRaoOM4TSRMghx6jPxM4T2lJTdu5PKgIUGhXkJAH8BuwPUm/TAFiLAjGU8HlLaIWMgOCO1Tc
y1FK7+Bo3QTPlSRfhWHjvZJC4TakNEsYUhdbZr8qENleBbwij62dQgYmmokrAhn7qY6trDVBeHL5
NDHbK6BSOcc7rfdCrlJm5pS/7xJ5SCIiw4UhrvZRHrPKnq1Jv2gUi+IyTr26vxkNJis7I8I32FbL
9dsrss98TwGwVpv97mW4HinIaYpo7XLIcd8QnjH6glDjH/6bjms/eO+m/3kV/vfIGW6pRnaCD9vC
yNFIqP2v+l3GcrbvjTa0jw3gfxkXOi+DVJ+rxoXW19YyKyct/Ll2bmLFOpbF+ww7oyRKq6NWY+Ly
bemw3SikMMYJ/BMjgGD6qQrHLuSlELeoBBXgElMuY9fEPsrx0HnQ4Dp1wnGx9mGZNddWqKTsQif3
1amkWMYVYOe1rtUmIOKO8HmH+d9c/yS6yB8vR5GH1QZGV0/1vOQBdI2CiZUQEhrCtHYK40VqjXT7
YaElRV0Ib2i46Om2npB2hZjnlFA/zn/kJozQE+zKMp5AeMo6FokQ2Q9IAYI5HuVRpHjjjhegtpa3
2XXzt+certpJgpBJP+OU2Ur9wZt5tTBcFroujLb3ev35B7JPcS/U4p23fxiupc4/0eLAX3TVE8Xu
iLSB52p8zJj8zuH7doWuX1VgcAT6FLsE+MhCbm6UavzRysQ6TzqBKt8kGUZqaFyHCLQh2WqgW8jZ
idS9mtfCfpyg6/rRmBPFgRXxFUXpKHGmhj+bx/n4ybkli0lKTu34sDr6L5W8Uwin0ClbXKjic+n4
dGswtkIiT71lNy4hrrg46shZV8b+eW4eT+mDo1kD0gbstLsCmQBgC0PKn/+B7D65BfB63kPTvw3G
lrHIk0S1XGIiGB/AAKVZ52kKGOxaOFVWmapATSOTstMW4s/jZHzS0H9Jrarpp2n6OrO/rJreAP8L
18VQLQ7ONqaFCwH/IRNbpTH9ejKh4neZ/IwPDNt+qB6lSTgpJ/M/RPpYTJ8Wl6pso2sSWtzWKKks
+x4SgP5k6qoQPKNK+YrX7an82aiYZnQaDl1Jk95h3oyWpk6eMTJHJSJBDgytUvNc/67jAmD4k+P8
5r9xScWppySUiSN79fYtH33i8VFnH7g091ReudjVs6bouIqkhkBFSe+dkcwLEhp3MIK30kqmDSLH
n2XbC1BuFliqn6utb3nsp9hdGMdSpRn7dt/YfqyOcUNrGemM35QMgINhPj7dPCwYwE9+DpV/kh5A
kF7i3aLh8ev0ezv9I6P7iv/4YE50FOctGOO/P/ZoBVjoQizk9lRHtnzcymj4nytF89PwH0lHBwSq
mSoIssBufY0/UxTqw9jK54icFNvzHgQSK/O4qT8PiIPxxw0j13ksJdbHVHNVLGozhVMNf+xWPy36
PA3GkujrSAbaEpYY72/nVViZuea24dBozhbyEPTyhSh6Tc2ExCWqwcJ80Xs+wVWXfiCSkrxhfGbO
c213MHihHOxKnYzm/aMVFPdQU6WaJnd2Fxt6pcsltjwZYrfdgIBYM47P1Dv7i2nSSDxaCwGB7jb/
LyH4/QwAck3WcXj2Cd8S4r99nEgaGyg47kFjT/9Zdam++iTcAZK5rRG8APK3cPFlPXXhpSwA4qIE
gDafAkVaJ34GOz9ySZEvTqZc68ZsY+CljP4iM5oQIVFCziCvZATDIC4ev/8GGPj0qC65si3CxSH5
MZRYHYQ7rMChigzlIxDYo1nymtq3v/FPex708n9ZM+tbH9oMZNNnPPPA7IireZTjhqPVRNiArXGr
qe05jpnaEZ5gaLa/6GVm7hNKVIpbWAtfQJrSH8ZrqoatISp+e4Hj8cyuifRsh5kDFnwkQkDjNfMN
fbH7Oj7SFS069S3aQnu7mBCj4ZuGDJ+LZ6V7nTio+KzpjS6Cgmy4FSNXimpoZ3wJHI6Fx623RJ5Q
VnBPix0Uu6dDpZ1RtapH+saiMXZFo7cYHrPF4KFuB7Of6YuHPuO+Hp2XNuJFi8RBXwcJq8FvLR22
6ymHqo/jWiZTWUuDaX3pJgF1twjkE0Kr3wKMAyUmhgr0Ouku9y3uOvl4PYGQEbRp3mB4lD3jnpeT
kqpO1uSGBhAr2uMqAbhRqpkStglWrI7yVzAwm14OKWUAUOfJRVAafQ6bYhoDqXlUqwfJ8Ts24Lwa
zJwsgS8OhCjF9sOaX0Qrx+LL2LlvzjHN/QTSQvoMWkLpATWkVzWcqPRiYlIFJghLQvGb1hSnG1Zd
aiTZf16CEsWlwfkO3i7kpntAlURRAgkyBg6RJqYDpafSwckKVTfnqG9LbPW9dJXV0mdnluZriyP4
fkmwBYSru+S0zxR2oPT9LUxdB95uNjZARWyWlFEn0UIcNyiEQsaBnc06qFmOidTc7eDU1JLw2HeD
Gra3++qmVV5A+s+bKoDIRb3t0w52n0p3XtUqbcA9VxunftT4l81zOg721p0LtB9qlcIv8GyXrpaH
msugXhmQ8r4WncNjnnqYtSLQ6DpjNMTqXPzlKMQ7QssW252N1bxpftdqNsqKraQKe/ZwI3omLxwR
jr/tfRPGEujMYHKQslkXkkLxGeSnHUO4zkiAORoNZJhtMf9OkJF2NkT5lbR6S7bzB9/ui2dgQOWi
90/Aizk50x6OzxE4r+Blq+WMpZ19jKe6l/4pJ7iyPPnDOSaNunqrN7tYaEksMwcwQGS8cYw+OLMS
HJ2dGYVKxTWVrZfUyhiDD06X5RURRzN4LYzIa3ttux65FKjEbXsSzcIKHFa8y3cRI/M8vnN3Dgo+
hZRQtLA0zz4VAq5LAqDRmim7cvA402vvcI4HSO+iyJAZLgWuuf4GbvuGvvyDhyspqx3cRUqetu4B
BnDfyjxdLwicgYp85hIH0fPkaDc8kFGqA8724xz+NfhZEChvEA77Cvc02mYPusmD7NHGAFYw4x2q
1GoxaapLww4olyb/sW/JfEpjcxv12IfycfbedlQLdhIcGQnc4y7cJxfqpgAstciJkkEC9aXikymU
Hyvpx/Ns4hNdVjQo3MT8Qt01vuEdQbXw9+HqvJDzgT/1tm6yP6Jt6oElfFu50Uiv1pHnRPBmZN6i
9cPdn5N9Cxxs5X6YcAVAvX3n+3b870AZDl9KoKc+pi+0UgR1Ys2wR6cRVUFln6HYa8xVLXXKJtUZ
JaWfq+MureV0vjtRpeEqeFajJaZH0bqydz03k1V8QZ0I2+Q9nafc11j2BMNGTt5b1z4Jm3WKFLJk
FUxvVvI/vBBCJajlK3C9KD40zz7hlmwVRy7Yanj2HEY4NShqQ7pQsatrmowZC+9MjyiU4gPcIH4q
tNlLoend71pqZmBlDW045rfyWvsilMGfODarGuOLQIGBoKrOu5RnsT/d9WVWxucaBOQ/dF/CxNZn
QiDI9K1QyeRBuri9jkugVstSG04/hJk+rZODO5JiZUFwOX7Y3U4W0QSEhBE11f61HdZvSBXp+jdi
HXvHlRAqXmAFn0QN0gWyReDRQ/Isg74jTBxUiDZJhaZkeGyfpijC5yFK5XrQ/XiX4gjl6y0Mu5nz
Ht427BR07/vx9obttQGFk/JNAvTiGhzR4woBhbBBRagz45ZMWI8o43gzJDf+xypJTg6By+j303Mo
wJsdExVBLAR/dFZ9gjmj2uTYU03jj4dPRwBT7GlBivp7CmV9ceE07QWUEv4f67C4DD94vdY790Ro
cl3SplEP1H/AHrV/Crm14NI9oQszNB1cCTk93tOUpqtCaBAIrjdK5xH2HwpwjYjmpdwalFFxuIeP
fWJuMugbnPwuErbzfW25eue95v0yIkh864u/iS4rK9gYbXM0Ku+tC6rK6DHHN643L4qQ0wBJCCG2
AfUASflhVYsF4OMnQ1N4CU43PuYgoXN/uDjSEO0ZJsX1+Lcs1jSymHfolyXUixJEYf0N/9M0BRUV
m2fAtpttr371yDJ2Uhx9nzy82rBgPo1+BnZKyWRev+6LvuaIh82lewendotGwNYRqG9P11x/CBdB
no6MCK/bd4x3B3m6Qc76Nnivvs6TUTHfJ0AI0CeHGV++hwiWz+p2gGeX5SNZ8BADwsgMv9xO1I0C
iEiZq74T0gOlLRH3TZTcIFolaK4zB0rLQ/rR3nTOXrmawT6SyrMMlHKENiTf0MwQjL2+6DTpWOTX
9eeHn4FcLfuU8g1BCgqTkBhMBwfip5HhmivbWvL3s6vhj6p31huKiXIMXtgbVSkH6lixHBWaer0i
Y09X4FPVASeRrWRHWoWObwFB0c2J3e+tBYSFxHP2q1c0TU2CmfOgAm0NVxbivU4rdxWpxTPRpjmc
a3HlifRSCX61fjZA3uxkED2z5ClN6Nr3Iki+Gu/wgz8rLuYThrG9yAEDarCgbTak8pZhVgHdfQpp
IcCvM1vpTwJuZkwRUdQzm+rlB491xPKI+WNIoZIXyLZgnkRTidIaebYf2xfSDhu3calQzutAi2dH
BpX9g1KZ0klfTNQEHSAV9edTwYDHwk24XRSV44KAlnHD5dznm9hjbB43129l3XDrMMGnvkv8Q8AA
nasG74XK11/exUxKWvDyB8NVwtaRP1inUwiKowc2fibiGz3Yk2HxvPwFoF0Ys+ygNop+Dc2jZ1E+
iGWqbNZVRD9HfGgilapaTZyCOyU3DagODzgF2edbbz7c8elGbfuVY3+4ZyrZFC2nyNCMCmVhHecB
R5r39R3DNj5lGoImp9Tj1WMwMiLotrHObryWOAVRrjxGyQwqrBJ4znmxGxgPcDoGRDrmGfV/RX14
C71cXXh5xqPSgsqBP014arhH9dccrjQFkdsWNdh50EqBiihznvOuMD8BhrNdqy5DNYT3DgEGMroY
iVvEYcObDwbG2cLDTeG/k0DB4GigINcoTso2gPpo2l2YQqLmvxZypuPqvqQeh6OLhyqe3GsTOZuK
lRHphpYIY1tpjPNDxXzUD05rtnOp4+LBWZxOoczkUmDRXrC6yvt6SD11MAmRtexNNMpBJvV/nNyX
5o8R/bknwWU+cXi3/bDs8Z4zeIIJZlOekWvs8LUToSvcpNO8pJ/BxPR4k+YDj+eh4bQ1/p9dzHVj
MCn6zfbMZc2ORuUnMLyk6ds2WOfMp5ZJzBEgNnIRdJV89eRH9mL9NyNw/8MRjMlph3wRz2tq0PE6
5228LYJ91WN0s6XxfxMVcUvMGNMOlX2yr3scpllWcaoTyls+YX8Cyjbb6+o3UNECeCSHFz2wcoXv
4gNMxMjt99mSkxwGN3B4DxHYiUAHlzMnuoAAUsrc7MCX9o8NdySZ/R0oJIdAsMOo/zCXNbVsaBEv
StecMVYO+OkJqHe1zPDrKYDC1eXqoZ2PSPApjgVS5Fjc3UaatODb7v7MhjMc6eBbuZvCzQ+qHK16
UGqLx5prECm/Iff8mqHygTK/Au7kqXGXGEsRb6pbN+Ge57tFbyiuszx+bUym0X589eGimykTapBm
ZjtMii1uuqZQn8rLMX5lXvRtZ+d2s827X++4aowOYNBKrkIOiOdJtrTHF5+yg+KFO0nECL/rkYlC
oB71hN+xoWGzuVkrrSbxWqJa3GFxj+ASn/AuSvPz2KYb7WqeOgD1Jcc4/6KkgWlOCXwWDtmepZ3D
Gz5RmKRtpXTDvk9o5qJkfZcdxoOKTQWDb7VzONo/9fKIS4Oe+ZMGFlGZyTjUguAZp2QRCXV9RqcX
LgZQwSZmtZRh1MP5pWJ9vJbHDMjCxgPxFvS7ekn3ShfNzvn5OThwgdaM2FPFSLA8ovNeIla7nb/B
ZTU5MNInrdl1QLtTHZ5fdk6vo8XY4ZJSynEqDwphNxptuC5zX5BpLCD4L/DjeTRgIQxb3iwmujqC
9HU1HT2v8BR38Y5DLLE1Uqa7vT9qNIoEtgmzVsX69nzqTcW+fgQRYmYMrsLU3eccaMjapn2B/zC4
knkr0NzN781+oEqiwgnIBukOuqh5zLHwaP+rMMa7Ds6cUNWNMi5zOsJ7+ktLSzTacet5W+JtQORG
mhyFjrdCai5qC+POHWKmnppMDG+95DHscQK8MzJi9SAPLLUHKAc6cCWKf4Td5xKhsT66QgF76rgl
CLl0F1BUdJ/PmIy4vorsDGnIkLdxP6Hu2jxCM+keQEaXBopZIYYA4EqHoA1gAjE72HkE9KcQ/bR+
8sTxr/ohzEYgYjZ26rOCHwVMhHCSUCnDxWRj5sSB49NgtbEaP+u4jFDd6PCe0MogUGHydOHPZTQD
BHdkKjEFC02bWF33KqkFZIUWklfyCLkycD91Eagp7178MydDLoBb71WktTQFGLGn3xVhHjP2YwSK
5OcFUqWd1KvnIxhDUPNOX62S+CGnQDDHqfWc/U/Djg22DRTJPDSO45CAiLt5etYGfk1RcA+W5GAG
lELUdDctv4dAOU7TiD+eq6oojdVxvLkYPhGs31yGbsBdQLkMxTyjtajA/qaogspE2r4q5yK2UBd3
RGHi5FYdqXmMPJBOTwLk+b1BgbvKs3pa4EdqHz76eR6TIAystbWSwAAnmetUA9S4Ar7FDr7A2q4F
RT0y5B01mVNlQ6Sy3lp4cGbdoM/u5D8RKMl3JdmdD17qMq5CKtVJKc2rt/BBpXvIAyDI/fSitv11
LY1E5zZ87PRzF0hxrKdOxMbOtquwaPlOIBrtbsLLo3gHRoBNqScnVs8NfbM2OoQQ2LLJTZKGCw1y
jPsZy8BuZqVG6J5zabaANoG9lm6WnIGatWI6c4LhlAUk084NBRlB816lU2khcepBTfVWbHQO/PCB
tiNRwwT0zBaEJx3tgYDblm132gPdBvQctkj0fVLyv1JY8xHMJMn5l7Pf6P4i9u81svLE5b6KE+a/
/sipwmty2IqTSXK9P+KCjdAYJrMwhLZu4aGaloHWQ2CwKMI7OnqveQDaXZ0XhUcr5A1DmKonzT87
nXYjnXxZGCaIhzHviVM9yx3QNz6XnWuddXD+ukGPuKYna6zS2P7amwn+KVCoolPfA27sBOx+QTtG
mVN9bkcKUbMnkCE0rj6AJ4/w28kzTcO3MTOZBMrMPas8Ugg9JRMmEBon2Sx/nwkwoSIRtqnloatt
QQZjqtKsVvyyxHzuq8kVlLetm6V9Zcc7nfuipAi7sVc6gFGnMihhdlyodICFybt6ZBwDnQ9CVc00
Y7RMLaFbmyJhjXfrnpaNTqaXRK6r55IYxJ2Wpumvmpz8zdQWB2tGnY2hSOBBQ0MJDpnJtsWVu+ye
+PF4GZeGtS68xDI0JgeJJX6qX7pdpiLpbC4vZb7HJ6fgV3IYnbmVKmG6FbxHUk8G7kMHPX4R7etZ
/AbXrR9Hmfhb1b+4ZNCVV18jyzNINnmNZM1TvIvTyAT5BxzV9G2ZTwKcmsAJIQz67EZ+R/eni4RC
7+VO6VGxToJmGAAd/vLRoxhi5tMmlyyDCckP3G4frS4iQJZw6j9EMslpmOU7ANuMjST8GSRKdDds
gJEqOdNK2uR77XoIgaio/eE/B776nwf95Ax0PPlAWFI87ENbeoqnkXcmWHZsB38QwSaANtTDm9eW
3EKTBrhohK15L2+JJ5rCAROF/fucRw1UQWTQDx29l+Tu/RB9bRuO7/nKv1Bkv9FZoPXqbARH3SYd
awUuMwSWW1FBCdx3uSfd2X20tpb0ZcU2zKysjOGuEeWkU/C1zqVFZT3H9ntm+VPuNUsJsN608cwK
Kf1gWru8o3+syhXfVpM2S4xQIvxwZfyteo80aMPyue2H6LCiwAij3da7Ltv8p9u7t20/kAKY39oM
TruRm5x4OrJPEDYoHfStasjyR4Kd2LfS+wDX51LepC82sawn8Di7dkT2G+cMnUucblewRB1RFZ11
nNZbMQqn7CEHH650/+rpbcqVlg0+aAZBbpEfX5Euo8LNyyXomuQdVfpsxz4xRivkjx8WFVbsU7gZ
G8t3UsdrP+Sv5mQg0bCUBCsyiiTpnCgAYX5cs+tB49iUj8GzvBAY04NO5PjsTLdm+WR72pgLjI0t
hV37HY7cjSDvPO/SgwD/tCB3gxlYIhiiIqqEr0WM7FGKAb0tu51Japdw3jl5YJ7SjBb3vGpaapei
yYjdehOtarryLFYObDAta3hqkNmOYeKqaDi5/jGkNuONtByz5GZ6KA5C2sdnEmM0QokxchSzv0wR
Z8MuogDgNtk/WUeNDG/dTcQhnx3D+Xdt2hb8DFC1Y758qwcfIYXFepDpBlgmq7Ap+22BnOOgSmP0
WYTj6Mc4CMOVmCchYsGJ1gfaa9SMiaYzXdNQS0Lz0FIaBU4vlUt5853Wr3IaYG6o8WbTEMQXrhj2
msQhKrNpgtHpUOSuwNi0j1HzvIRrTiqD0mxo5r1sdQgiFjQN727IGQ/l5lft0Ow2xSRs2A2wzVT2
8wdcBPIuOYt355RWheSENH9JUo1YkruMlpj0ZKv2kyeQkPrFRjQyhyvbPQgyYeZmDCuhYV3d0Y3m
5Kd6SH5To5W8qsyfuts7KRTbV6O7BPqdLUSy4e+aRrEALrEXXZUU6V0JSvg2aFvoBu7omPoIpBt8
2IRM8jig2jU5/QMweCLioDnezVC8ukivGjoIIRus60Rh+xwQR7uO2mRrCR8GsXjC6F2/FNPtbwiW
qP37Kq22Wp09VIGQxaABxd+I1nLY/yMr+8DkTsgOisdwb4j+cisNQusPSe09xzFJgYEs7nzuDWKm
Rmvs0+V27iwvL0Pe8jJYQsUnnSEIU54eJagchcQrmsVWVxYs+OX4L2/7nzReowhnEcm/XQ1IVIXd
H7e3OMZTrl1BqXBU6Zxm95ROCXlWKE/yMqnjzIruO1gNkeW5aL9d7i29zYixugQnTE5nQHwRRfEz
ZJfcczLVc4PCATya/CJjUJ/Cgr18VM4jk89Q2wEvZhKK10VzoK7V36fpqjet0QTgeWwGXtZ2LRzW
qCHYbZp0mxH/HR37rj8XHUmZVL+qLguTs/ueOpygINIV4m09BMzkhSnfBicr0dw0ClsfXBm2Lc3a
ayNskQT9WZk/VLaQz9hJM7Cq+wXJzehZsYaqCu5+uROqkSuoaIIQJM11KeQDwfN99SGfNqzFytGI
ose1kIShiGq/r0LJq0Rzm6/kzEgkObwaFuVTYCIPLJS2Bczw7d+HEBk/nq5z7TBv5U1gjSMSBd3u
s/pWH5Ake2+L1XqOzKzIN0hT+TtzJZfUmvks8KpfkXHPlRpJlWQhRot42ezOUwzaY2GgCd/BLj31
MM4PjQF7SuE6NxPPloE6ERSFGBkxoRlAdx+vmlsEzI8Bn4dgR4/2CnHKC3gcTGxr+zhhBWp74RWF
myz3cZ5qXudua1zTq4KFy76A955OjSm4Sz3epwXEbDkuFz5qQH9n6oJxMnfkbcGhWwFs6J9tDhAj
ulcF4Z7aLv7/WgafyxxyF9GGOARlDa2LftBfzPbiDvFG85zH59FlJ5itm5qU+fAO7AMSoL7oBt35
yj3LzbrnsxewV7WTc2g3WlHWinnshUdkk9ABja63lEbX5r94HfYBtTqZzXQMU2CAzqXYJAhhmLgZ
plkMK72o4Xq/IhP9Y2/9pZ0tKpixlekHJGtA3I4fvoBkYlJntfbpyU5yNo9EiIARhEYv1EVye7wt
x+5lmT7ObVKq4h67bagNrrHVi2SbbAVKtZ+A25iDpSFD2iVG0MI19NIpERiOR9LWM24ETswa0p5p
e6pHWEhLnyXmTJWPGfymKVwcIIFG1s6Zox29bWx8lnf2uJXbq3lsOSW4AAAy49BIFFqsLSx5SroL
wJySewTkHbk4NkdzGj4Pj6oMlhIEQ2Ql3n3wzAgAMbTUWkwmLSjoFJ2hyXiUDMvezihB13MGr+gs
NYENAiGx8WGlPoM2QWHKwuJI4khePgQzUZ6oh/J9lTf/rTzdX3e4c6tPD8CbY+c0x8AA5jY74xlX
K5k0DhjmDOU0P3DlPaYIoSzHT5P/LgzKQER5n4Fbq+/uhRsVWu0Z4cqvrSQsl6r5OOOAgPzorvtH
vIo4UjMwvxL/wK1pLs03+xhTMT9Ay2eCZm1jbJWWltr/+6oKsTf8QtZiOeb79a8hPLTbh5ucuL75
E6eHB4TtaIYwnQ0d25HCa3YFitu1AQCi7jbtnGhz6y4iocdqBdC1VagE5ZjYNH5c8Jxb6FDQRCr7
fKss6RdklLNjgY9WEgrQ9TtRIvFNUMYXzaeBWz3S+U/Ct4bGO/Q/o7AUMgH2mtLuNM3mvSAiuVY4
9lyeHhSdpWq+k1ilE/x3hlNDMNbEoThydZhHk8+A/GOaJffxgDSw7+WYckOqiiR6g7NitzWA2Nl/
8rR6L9PEzksr++RcQmYqkEU0ntjD0APDxehtAjdKTaf0E6Mh3H1S5s0SmK26+1WRRhqiQ3Ifuqrc
DhdDdQAJ0DVi10HN4BOgEA+hTK+Onpnu0F31Gsp3CG5SLACoaf+XQcJx25w/XwRNGxSC3ZG7umV4
hK3A2WCSPbF+JJQra/2o95zlyMT7XTXDwCmYtJgNAT1EB1Pp1GtKXWQHP6HpgikTTvWuvRjdU1qW
RpUHUV4TKPW6fW7YuVD5Nzqqo+eYz4cmMTLMvuva9E9LQirni7+A4jpMkw3BhS/9taULzbcuPeVH
ks/TscnIj/0vLm5p3Rsl7lgRnYtP9vA4/5kazSXd3jqZK1v31fNihqDF3HpBIfhse2+4I/xwcgMB
8SpDwmN0iHocUyfVHx/gyDSmkHyWW++HQhfhWejmwfQsXokNF6qhPO8HaQr17S/8cBUeox1+4u5o
hJd/BA9VybyGlyJ4kZ5k95OTjX+gL0QgUo3KNeXkzXpKwf80eQ6uTANbIBQOMo6MBBdSeITSfzMH
Yeuhs2gSq5Ohdf2AHMTh3Wp99FoMCf9Evn7iUQy+sXwCbyOKhtwDp43Pia5GfARFU+2XIJf35RL4
jHVJurCSZyOO7fAQdWbx6ELKoyEXrCOWRZaMfXFkxbwDLk6QhcG7CrOGRh86sabvpd4lsgls6/nf
DZckgqWfc8Li4T/egONOgnYatjEhMUCK/KQPyLnnlD4YzOYMkoBbsetoqMa4eomLCyM0/dY2mCL/
RpvjR3cRbXrW2HN7VEWH25c4ih4Rrk223lkFWLKkw+Dn0fjWotrq9O6xcCDe3wpXfHizx2raOhU+
DrB774FigZZXgJ+0O9D+EQQQrPc15mATqV37JjdlYGrcTQg7mEnM8hnDSZ5B9k+U3bQ2pzeUYlSc
31JWfOOVyjmZZJsPTWQU68kxlG5yuY4QbGs+sc/t6IOWq5T8XuVnBojAP8M330MJt7+6VVPTFn0j
wRz2XcbHKCQjpW4IY6kjMA9JLoP9RCkIOxhaxWleX4spm5SCKKFZ3LULzFVoH0PwFmcEEtSSA0R8
LGGktgjE/lr1rlOfA38SzPQIMO7OO1aMavhHr6jFzw1l7LURICWU2fdlxTmWQYKH8lxUI3iBgcPX
kBf6NpZ1lnbHNZtQIhOv8P45IrDtE40qkC5NwWaYLmgCYdLg0uPw0LbTSh2k9gQBxUf/sKfeeDW/
QDgS2fmg1/LNyO/Y6jpR+Jjb40OcSfVbaHBJJe3LbuitWLDJQ1iefG7QDrUdxNmaR+5Q0baRfDRo
LmsSXC9C2xs4zEtWIT0HYu98cjZMpEwq0eRhlxcscrEpiYcfwmxLAFB6NOqQMmhZjEZrYhavaIai
SzQwPtGLo634muDMERiR7GfKMMlp426oCRmhv5KzhpykWdf1heuAm5zy0OxyCt6CuMl9eB7F9F2g
eCVNCVKxYWrssRal8RVcpoFy9Oa3bFJHQcwYe7fo76md2yB6W3IeDqzkCMzTt3Swkec3wzr5NHtZ
HAwp6tor7grVUH8SxjD1p1Gz9R1dDyzUUcnAjwfHJNrwSrBc5sEcFxUGOFV20B+M+/0Hc/1E0TfD
7WpPznhCKGn4XWPYrk0xZx1EsYQmvqbn+f0Gv8cRwyyJ3wFSUJcmjWcrJ6elbnajbgDvoJcMTr20
PQg7uToyCj7d+euXDjxwdnKa2uxOi/SWBV9EN2Kr5NlXjnWL4c7V1KE8kfl4thUOvgQHdavhbP79
ctyD2OaNzynTi1Us594UmZZa9JXwwPU3rLvRSdsR30ZOGckq6kfUgxpFtAshvXiOrTHWmc4qp/GC
Ffvi3f7RruyuMuhrxKxWlcEY4G/0sGOBmfCO7sczz1UNAkBsWpVhr2HtTg4hjY/cVLH2c0LbqVEN
ZA6qG5wMzXoM0u8zVwO7KwQQgYDbatpFdrLVMRmvrA4Fj09MytfsXz7Amakd6kTKCSG+dXhPqbCj
CiMHLOP5sAmRFvDmlI+/zOAu9fRMCUI//ExtJQHPUQcUdvKuWf1Gs5xHk4p2AditlzLCl6yDEKUJ
W912xla6gy5jkDyccD0CrqvHasjxw/kMeX8fRILw3hEgUQsuw5J7Mwi7JXESCtRwbdlNKSFcEEUO
5P61qtL3T/hx0Qh+b3yIqaqgJ7GgELRWFNHdK3cd9qyfVD5RvaHYDnwsVJj2DmSJoh6oL/2gs3Gh
0/jn/xHyqnIry0zMk76ZPAdFRdVO2cTXTj8lhgYmoLu0sKjy2tyeRwm2d9mJF/OvttJimvf2rzDM
UKGRSJsGFc2MC1dWPcicQ7/Pb9Ehyjn3PjDQlWZ8p5YNirJmqwFSwT8MF1F6lvLtD0Vj9rCKPEso
jUw58hUlYhkYnjoNDwX4vBSQfiLyMtI+JuZ0BWxRhZUbRjLzWirCI0/yk7OxyMZeGTFEMDqZ5FI0
ukT02W3V3Lwu3XtyA8UaejMBZ3d6IP5kezZQwKOvP5Tp9ZgyBo4C7BROib7NerNMlZOnesS7jVhV
YvURuCH0ZUe3GG/aK3Tf84Yvv3kLePHEPRcw3ysQrloNp5nz5N0otxz6x1eQxkyeLsAKZbPDunkB
WIZkv4PO9xz0+Y86DcIirPnnilactmJANHqp/9q8FxPYQLQpJdXczLm6EH50pCualgB/YtQQE5Ep
P4cCvJVZjoPF9WvwA0kuzkwLas3/EPJT/sZPnGKBdMM4IkFsat38Bx8XDFtlZDL8UyiNjuwl3C4M
6XHL3kTrpjOWtCHVhoopwFO/bXIRU28gHKaqKVvbpeOLsOhNTObQ9iJ3sLofk8kJzxB5KF/URtGf
x9e8PDp9hRk48ab+3tdXU1G2ddRJQWNAryiTACJotrxC9iVQPfwUI6lZsgHa4OTLqxtC6cpZPctn
IOMe0ZQzlWu+kzzW4dyySB2lsc0LgEt05Us0Fjg7eXtAd73Ra9NO4M9ot0ZF7vUtzFH7F7c+wS9N
vOfm57Zq7DipJQIVimQxHg7Zu+paS1bDV5DZHmDS1Ht6ISyOCXsXAqYh0s1lzsY5dTMXboJoZ+MX
CNAuinn1E75iFxN+u5Z0+P+BTifmzj8tRAnKEu/b+kgLIlHfOS4RVAKjDphyIcuqLY5LqxZBa5MD
NQDrDiiw3zp1lXq6HF/C1kOuIidb+meAGlrUjiIF3h6VEc5zyi/+V5BoCml8QUxGQhVptYs+mfp8
iafokpSH/pDTbWF4sz/t+v6KJygmtasstuWkRsYIk3/3wbanvQwPNMNQrfupXPjRn+QaJC7vEEyC
O36wnwpumsMBlQmMV22SqRPFh4R2vo1ispj9YFQcbuYKiJe87+siQiJU9bORSv2Ih6T4RytIvoSW
A8FgqhmMsDweeJXDDJT4waXoorQ4Y8wLFn3q/tdanNubZ68oZJS5xesVZNC9hTxP9RC1eS09OUw9
d3cKvBP5jFpUrK5SYYz9UzOfYsVpi6XfYDFXA7VrTdzjg9PzClIpFJxacbKec47cs0EJGRrMFY17
UxqaqQSMVHvhsK2BgO1pEvPMiMZcRoLjkSGDc4c53Eze9vYZELUW5I+8onjtPe5Oep+NuZz5pQ/W
kMjsaxQDd/3mWPs/g1HFXc/cAyTCWZad+Vj7zqVm/WkyAR19BzJJJBw7BPadp3RysDVEHGIzK/eQ
HnTIiqhzfnM9i0ZcwRci6JGW/a0bV61A4PFIY/jOYrutR4mDAPvWSG1kpjvgZl2Mk+SKPuSlLSmS
YbO8n144UURzDw37bybPmS9ZdiQBeLiqs+ubLabp5JmBIJ6oL8luBBkGGhi3/pcDqmdaDLGcGmxJ
k/Qec5TqF/yhQCB1lKlZgILL8XUVJYYVufqkAFCrthA4ZLbKYLBDGASBD+sTHGzM4GS5Z2Vd7L4+
QJI2PEN9NIFQaNtaKpMD39xd4ZIJp3iZnKcMrT3i2RyIaeQllXPO/xsdLeL+V1rj2wyAfsQAvfkD
FcVtrfdizEP5P0N+Ch67USRaCMZUqE9rilDpZsNxvgIPdPLBYOm774Zw5WLoTgANzt2aQYLo7fO0
OsVGCwOgHWoXHF2KTgSpMlVAUiHOpdWaqXLEnOh4xgXh3B/Acu4CWe0i31ivteRmMGrNhPAf9gL3
mvwDNqErcoB/yT/i2TN0N70Y4nsvvD+Tf1fx3zxljvNfyUwp9kfgLHCGMQUa55NOJ13ePx47axk6
qbpL8ZyXAwwZLeeyDe1SjkWUl7h89FzIoldBW2Y5agF8wDasBp4HcxOnIBWypNjWabotObjNaE0P
BgWRoo9pYXS7Phsp+1vXcGla9rehkzkoeCKOujzgMNIBlYCebOfIevoHvb2ZBCGRCgTgnDHZ9dvI
TxTSXnlRmfq9mnp9xcGBUL1jUvN9iq9z0sMuXsYdzAB5nJw/2Ef7wbfO01xcfSvTke+Ll+BW3oUe
ajaBb6HN9wVJGVcMhtM8STszgiWEjs1a4s3A3taYZGTS8wNJgigY41bWWVr+mS/quxdVTVd97nvB
jti3QFJ9dzl1qhP604tomjzR7QXSL1gML99w7RxTibIktZP5fV6/yy7FKVw55Lx/0p1+NoR82MXO
fD+lct0V/4oZzycPnSPIpI/7ExdknHwCg+gfAcIHGhM/9Lnu6jASCmUdF/Vw2TIOvXgjPkhYSsUE
4VBsFr74Y3zorWAQo4wVeeD2PuqDUtAo8IWoEq7IN49esQAqMdiUF/Mze55PJhjzbuj0Bypk+Uhp
fUbYDgCCogHKRG0WyhC1qZnl3PKvYfYGd8zL5OcT7QSfSq4vUuk+EZ0oM4mDk2U5NYqb4/Mc972m
786pXdWvcnQOoWjRXKwO+6XIeK3KU2IlJB7aDBWmj0mN1k1u5dqj3dUGAEyYC1z5oVlqeNs0dI4S
w71HdGWUzq09jhCkO0VxWrvMa5v8RuS7X1eHXDXqWhX0btsiEkKho/chJy3nn2uMBYsupshLL7KQ
f5BBhqKAMptpQTpdcq/KMIKSezioO9w4xWElJHTORd7r+k0J+48pL1pcZVhpPACAzA0B03JVe37S
eN/kK++IkUGlEAbK/AyIZUh4lCsbTnGmsPGElyy15HeVHp7z4IlAF6xlJbwexlG969O8qbLrslkb
3h+0MMX6TdQ3gmap8WSmRuc6GuzsXWCZAKefXhJAf6Thtd6pfcEJUCpdwATh5tMpx4/8qzMlpitx
9bkvQxXmHaZVPhfb5BRAnguE7wfk8dQezOrMRSAgOMz1ZtOicsqVL5KOeZwkdmLhwA3Jo4n6XTdF
d7H2FawmEMfysQlKR7lKx8LYsczeidTI1wXdKrGO+wE5DQaFcbfzNoyvWtqRLcbxWj0HZTl81PK/
NlepawfgGUbe8+8nkzEmn2ymzvhDEV9Q0tnttw20we0KQcF2o22vAB0bOWqNr52K1KVGZiU58jJ3
lHTYPzHlNvrLqxZe7CzqXAS53kM6hkOs4xOlq3f2UbfAehTlvfTj5Yn9BwYhiycTSyyHDNCWJxJq
FqcipM0gHuC9mYZTOJB+Jml5pyiESjGj0ZtWIQI25VVdYyvIWlcHQ2WoO0XuMxhNZ0IikOrbk6R7
96hPFsUIs381mjple/ZkkRhFBnfrxOzFRUhUfWuGEm6pbAXmxCwgeAbNhZWc3VBzZvDBEuJcow6l
56VZJvhPU3gVg6zhlqYQqyEgTf9U8Y445KLB5ldLzF3xTyBP72MrrLuITTd6Wm2iCGwbi4Iplgdk
Nh/BbLR0XAxo018jFq+yLeYOxIRTh+RNIfZChj1QMKNdH1E5CmM/w8dT4wk7jEUalmqEy+wZ5qZu
M+ga0tF/piFVm6htsFiabZfnz74bavxMiXXqpv+ZKCtbqJ+CHVRvWuXZGC1Tgrp39otQTcuxqGW4
lGDJuNjOdBZVq0DvO+wiOhWvAtGxEVaqPJCFXSUr8eWUh06GN90Z/7BMCJikMbzlOr3Hr7dcQFhV
bBeu/LnpIwIL1VKH4IITfelmKXO5k1RoeYxgDANKg1kkqOt5XDp7sJOOoiUCQOO7LH3BvMDTS7a7
6mOC67gdHGkSsL4+UQUbyMB0pUBtOBdEihhz06HTCCwT+bqF4xTBYCnsZdbXdZXfcaT98IyooF9a
pKC1/XvCo0p3xG/KFolFNw1XONhvnrBdkZCtkExjS6AI0Af8D7SAWY5okypQ350yJSrnYsNanxlx
di2wZtMdZS5FeptXQwUhezT1hy4O2dKuhUx6JzNBFXRjv/vnb7rEtYSfmto1TiACikg7/IVI92i3
rKMYCFPTl6Vv9IYhN+BuqcWnDYEgNJCa3X6OGickOQV4VdQxtc/pf+usuuTulmQdcR54YhlATWSC
hm+BwVmdUmEmnQGCNN1P2gOY7L+utWX1ADF+HBg6okOWu+V04luGmHnIf/6Jhb2+BHrQ9Avwyxo0
sSSSuiTnvqjd5mNlsgk36U96EdgN6PaBBAifn7+QSl4iNT+kQW6ezr6J9OXLo6nRnN4Zj1706ktt
vDSHJ67AmOUONl9nFrauyEd2PRsxObjqvan5dyg3QtRi/hFoXDBynVdWsEhSPqHGr70a7WsEPux7
RFrN679ve79SEtBeIR8zNlNeOWd8/n+Ry48UhS91e73gbAgs9UGX5IdOXmGDYujgf5IEpXqvugFU
VVHLaCP/7fy00cpSbGSvjv1dOxF1tN23N4zrdbykt1nRXLSia84DiArq4ol99AgLdAaVxn0iAP3A
NedMocGkyapKBmA0JziTdu8DMR730PqA4kpcBZRj8Sl/bZn3mpjVqE23YID0IWVJItO/KWQJN53x
DJZYpCoOttWh+couXLQL/x/nPJpFnBR1+FQsIphPMZkjvuMdpPYQ9j0hinzduTFEXybvjRQSorWM
LvfsSaOvL1Pz7eetuMSaKq8Th6f76Xeorrc0OllS+uAy2npe/y9sUJAlmczUbFf6tDVAqDipsZgo
yGm0bJ/8EY5myqG1P5+mcc5DpU9mVIp+o3E0uM4DyerPKgcp8yHQP0vv4hJyeZznShXTxDksc6oj
COuNqckI7lw+lpwkQErLe/TDIHkvD6u2IScd6PNey3XM6zXaBZzJ03fynT8oz4m7HhbEHxWpmtKZ
Qw8uGyXNG3ckHcfJK4g5pJHfWhdgV2vAVyQHhVPNoQp+ues1isZ6njNl2LCoqDMvashONYMkIiG+
4ixmISjGW3oc7/3jOvD+VQrUxGvavwVySn4SeuUjOJbw1oM1I1e+xUOGcLuQ0WtaIujmtri/fN4b
j7DpGQzLHuv15ZDPxeq0LcI+JCILV2U95s7oSTFTUEOUqQkeNxg54AhWx7TdxH75cwR54e1+i7DZ
QDkcVaMbCRPyEMbLtaFTXE496Sa3C/rJO/jO9pwvDBiLYNkHa08FH1j1B4i+B9s08dXWH2uPDvCV
rq04ZtVlpgHSxyf/9nBg2KntWENuSsVK2HRNuYE+5hFBhM9LkKRdBoc+OMQex+Oggr8/aOlfVqDk
aFgRPLE8dGMAwOKFVj2b+uoKGu8nCaHM6AlkXul7IFkbg9oK2fY6Eap760UpeBkKvE1qid5aj8e+
fQVfJZvdqVmZemoVvAXPssoteAeq6sl6JNmw20ExGhIV518HIaO2Kof5cbN49xDQs5JJRg3wLQaY
g6513kvFqp74UlvPAij7BRQpuJb3tYBqsKnxkNkdYr5UddVG1t5k7nCwGLhzDcwt+pTbS/nobACd
4HIAep0Ibvi/iy7c8f1uoA1HLsjRej3f9PHRRF5wu3thw/0OGj8MMlxBwQSwKco1sBJ94Gu4zMn2
FddaSlEqNgJHgrvfVoHgA2iLKzec/eYQPTcbCI4Uo7YfFj1p5dkw976Gnw3vAaN+o3MUplCLBAPu
4Uze3yuPenyU9w/eQyppWp1l79wR4o1+SlYlHSo9priTwGbyNDB0oAJ9Lpd9tS6yklZkJ/QCnudj
MtdR47nb+wDUnp62eo0Oxh5ArVbF44wXeNRrp20v50DAoQMUaBoz5Lx9gmeN0++PwtUXOa/j4MAX
6mLAPfB2x76QspgS2vxvo9AnKzbYg4yz7Fgke9eKSSthywRn889AP7mdKnZF0OU4+brBWFopsrP9
Rz4/Rvo4fAoEsmPDkRvl2hpvtWdOpoLGDqdqIDlRVd6QEWM7K0GWn/U9ucjkX0yqZhuz1Uuu7tka
Ao4FQauomeKQhga9jy/asE0XysOpYGbop5MRRTB/ihnXkq0pBBaS2BtAwM4xsC/sWip8iDEOVJvU
cc/9+AR6sza8D9T1EJWb05vxiDXZm89R602mWVr2XGyB6HJc5FMU6fuGkXi+qttujNrgMC6DwbP4
+tc++exIiOYH+nZFG7/fLZCBtHXBAGEKeDX8EVh6nkOF1zjitYcGVXs0DROj2uxBuyyh+bT/1xeW
Z3rBiLDLBCEl6XbJVST24W1FeXlFvKuZByNDwchsdyOAK/Tlo9UaO2COjT2WoKUaNZrvEB6Cw+1y
tcpxsAdtS5JisEwScWSEOhsmy6L+sMORaUcVr9Dq7LLFvnjIOwGMl8kd33hDEQBThD9da42qXRRZ
xWyi1E8MMbtnetZL3LNPx+B3PM68tMHcTYMpg/cr7ZhWEMVqCVITJNnUgzRoHNdI7HxvqkiNvVaz
TQmvJDG4h4t/OOycABDOYquX85+7Vu5raph3gwgEbjaZn2cgDOJiGgjav4Eh9ip3exUdasIaC/0T
V/6/BPQAlkzUzs2juo4LHQhtY1Z30TRy5IuA0TJg7C/fBZuNPyNhvpoui0roOgS27aJq6Cu2ol9q
0VIWybsYOwbIf65pWrFaX2U+cNn/1jxLcqKsU0v6y6+fJkb4v5m3mTwi5ugLuzxsTyH7LeGDwzH2
o7CFexgmFQB9k3swGDqNsUWf803uKunlTGmiS4iqu7UPtvD+5v7KXx2ax3oOZ3R9G+3NqSb31oEA
J3/6hkvP9TcBhO39IT76D9/KElXYFEbRNvSGmKjqzRSvK6OVlcuhWmPGTHP9gnHibiAGCMH22ybL
KrjZq1t/GjVzIah03pqeDDX9GLhAJ3SkGbJcvRYKdz/yr/EsmvYTmuqijfG0kRj5ZHKyL9FnUOwn
5G3WOu0tJZNSjikSnc/Fdusx3qOWBWw3pabVTmMAm+JD+hah1lR6YuvHenbXh97+K2pVw6q455NF
TZ+BE2GUrbhiMm92v3VcZbVYLfIsbHKSX+SVv9i3ZUv0MiMwbfO0WgkNGTo2cLAYgqMFXAdZvDai
wJe197wntySsp01+gYfqtkJxTHjXMHgrzqaFbbR5byZIlaAE01qhTrE6Ji4tlivsbzsIkVIopVZV
bwYpRaWAfKOqrEpV75Q+VpRhIurF2BQmcOPDER/5HFcS8tUUkk8djs/U6rh3sClhbJ+HsAnfc2F1
df/qSjYW+WofcVTU8wOsZuW4k5EKOzZLtQuxIeCqjnK969a6uX4h0evTPfAbf/nx8LRjlQE9+B5V
f7oxx5PzYiVA8gPvhNPLzKLqTfYRKFd0UZdd53sgg+LmD2UZV2Z3uE5Iwma3wQ+Pe5A16HI1wl53
obf59fEePcO/AbUhO09/IKysnkz/TspRk03AxdhVMoftQPFAhWnM7w/MT6C5kyJ7npQWeOlBZce1
dGzkTDPaGlStQNURha2yoYclG7W3PRxKDGzYgBIqS1XkcS0zwmQm+HCR/N0jKm81LBLS2qET3wjK
7fa2QWtBxMv1HmsDK+F5IRW0Iz24CmlhU+Zjxz/8joympHtphnELv6z3XUEFWNTJHQQvLqinolot
xZAWpLH7ThuwPJ5dt2sjwaIcpsafRCDLSEO3cEEDawTWOQMyefFAwC3U/xG5dzX88zfWXqeNUY0r
JEJhpgattHn2CFrNzYlmSGvmmaSkuxoPNU7sGIcrZK6i64y8/dxWDMFUH4k+RIIe6cR3EECuBCbL
i+SKWzImrY9XWVeZAQt6fTthOOKkG28KpI4GwdUAB0NYO6PhyGigfkutgF2pQYZfdUsPFbgkCsum
sWoIZk57R7KufKbIilRDdmwF55mJSFlEurTKl1hI8wNUHg0ZtHfKYvLYpwekKZNQd9/fxDXat6Ku
s5Uf9rmR2f/BfSlLAx9d+SN45Oc5rhM0c+5z95vWSxRQGOD8jZj+Rz0YRu47bb/FoZI6z6p8o88S
FjL1dZOZZc70Tiw7eyJqIb9KCBcAAAXM3RbQyT/ai79JOyDIqc5grrp+TUghweDcvr9z3IIIqv2u
CgzKyDJcBDJeWw5NQXRhOBQMCQH+MuokJiBotTrLIWbDAZfZvhoO2dSOzw8rD0W47bOjwF7rWTH2
X3rPqs+N6/Lz91CsI168ccJvIlPxPzl8Gch73JEBhbY+7k4fhVZEenPT0BABc+tuxJE6JZoYqppJ
fXhu2lcfqkG9A6j1Pexd0my5tyfOaauUOSPctvjFGyCWpUYL8SXvwRAWOWqkw023auuZL7Sxq02t
vzapW+EC5/vcHAAZwhct0gr4oaxWqJD7i87BIMb/0b6891hpFSQkAqY5h20a6rsz9lq7IHNU2QaP
7KxJderWYehwdkDH93f72P9yTgW3kP1yvczYNNokDwqU0Ti/75YN8ddIvMORHcFp/51MFQEfygYD
+23TjFveURv4gZCNjAIgB68m1A2Af3tL4+yPDRheLyZ0Q+h4MW4QBa72wFvrzoXc7AaX1qqL2eZ4
rZyzHUkT2wNot+enzujj2huRhBAMIkjmcCgus11+nuzxKZrXDIQZwT8fXprFZoG5WONnLTPDDrsm
mj/h3p0Nr4u52pRugT8tUsW/RHD0DUBPROFizXaK22VpO0PxibsK/a5Bv5eX/AnsWW7JLu6ozuYI
FMbbvoVeJ39vm7xSPMgi1g/TVNG7WT21txa/ClKCa2s5zmzU1aGn1ZnkEBYqOsr95B7O0FCtK7WQ
4HrQ7h5fJaPQkoyu1riesU5qakYz+jrq10Rk7YDxciP7RlEOCnskXTuw6g8QccaMAKeShii20Vpk
pfAvb4cCcDBOlGy6NSTCD8D734nryicRv+bx2KwrmegZcdIN6oKQYRGOjGLO+eh9VXvdcdM86ScJ
s1CWFxczZ/DskYOwxT5o4DxJZTH5HGR6iAhYaVMlmsJsz6YcwV2UIZzSdYlWIel8Lb+9CG9TDDCg
6pqKLFCl5+tB/uywMh23dTumK/Pz1nIaevsqTmP8yfnYBNTlscbxlllcDgl4su3f0ap/dYtHbtgc
APYTH6rBZ15WkZLIqWiU+HyQ2of2O29VYNSZiNezt+4FE6VWGuM4SqkPPv0g3VEEGBsTJmoNX7CP
dPn0Buv+x4WXelx7Kny9vtbB1uWTDzxxgRMZnC0QAk3g19P1Tq5DbKfzD32SR5VcQDlBWvQwjgzw
a7IyqVXSPcn3RadQzdJfRnT0NDmPWUQdeRJsVfV/5gOzOENnrM7xQq+5AilLB73VRA7oiNGOcQrd
q2HACxDZwfYGtjqxH54kZ8fG2xOB4K89rN0QuHnRPOudkVbR+ufnEV7QBXgr+kxSZV7avkQ+Y0Zx
e6GVOl4SmgNKtaXvrSe7OQlaansypKl/eapQ6UCUiUPkglPTxdVlH/isz9g+wba4OGr5X+W0/Z8U
v4CV9JrElbQmmtw4g+9eyTGPl1fLpgonwfAtE0lOOxWJLfkNWPExcsTVZ0t6aL0w8vKo2RuEQfjo
TlxsPb1Cvkpckhy9HeBowhZFbNU/nDFO75Z2NU5VHn7M96vE3k73kqX8ubwMK0XGDaZWVM9w27Fi
AFwuTHQfo83giCFG9QaZ/5VZ9SXBovouhFpkKpl3TPlIcmybG5yji0EFQ5B8LzcU0HpqL80Kz2S/
aIwkPhHFvrKy3F3oP64uN+3TFoAj0Jd2AO+Kp2qgIKx7wNZHKUiLUoLNGEh8/kPiaGTNnKbN94ri
BfqYZRbxXYeyI5035ISM/kOQ/El+WQrWbWe//gzKjwjaurTsrYWye/pUl723Dl2gQfMPnPRQaVBs
SKluoxmG9n+pRdFErIvTIGArr4zz0G5r1m+ZeSWG+LkB1XdfNb9B+8xIXa/xNwuwlJ96yhY0U3I6
+bXMGVPtai3+blSozjhbRtHvywg+ECqreX/XOAXBWH5BLcbgtf8Qa4wJQPy092fnrg4C8/uBLJdq
odqUTNz+J5XxU2nge7lPwGaC48D9F3iSI2CQQvR26mw+4b1phYvp71+cK8jzSotj/2lWI3yPc0JB
B0SkIQ4blpRvq740nZ0rswOa/e46gR4iJ/glEOyAgpMHWhasYTmlWZa9JsX+cU0Pj13PY/3Vu9NQ
3dNWnidxByu9pXLgtCLoCv1VD8I+3tQftccvow16YsOob6A5QjZWOtkvoteRrJg8d7Qnk6eBQnT7
us8vAR0TLhgweLSpQv7Sp2hO+hxVIko3UAD938r9qlWEwoH0L61CY0g/JuGFEF09W30i45x9wfBY
b4YhuIr0utJBM4XnxCQhxD2c430TrzYZDWRYD/04+JCurdBfzha4hLBklL1/bVtYy+6cGS8aztzP
/gOBv4mclQq7POt1zwi50rCLny3sSvmtyJ4b3RlNLRwl7rKv29/I5fNtLcv/Hf2yV6InXnosuWXe
JQ8jrtdl9xCNI8PxbNM220G0b9KzfF88LTQVXZdQDDP4FYO/Yj4mMV8Rc1wtWsbfzgvbn4OXCvBj
Ck7QEDBt8o18854bjn1xyMQ0HSoUMKqHF1txqBQguJBms7hICnuC8pEwcRzgeCHn+vsnWjWQ6sJj
ks6tcPA/xl7iTgiFjhi4044c/LxEGiJrWBGts9G76qRhbfBdbKWzxB2NCPa5giB/8mFQ2XwN/doN
tba2GdyQbyavxZNvnUsd5WQzLA8WtPC1ulVKnKjG8NDZOEunV/BBifK8yX5uOb9VQ1QpugJUArhm
CyE1hy0K9DxxoJCAQCFomC0PNrPXDNkWufIFLMyONi+kFwK5k6+MlgDkADaq+waHytWuT73b69eF
7c344R5jyScJ+oG9jRmYA6OC+5Cv3unBJYeanWUzHITOZAGKXKkQ0gU5/zbC3qaQw81kE8GzgPXY
LsWP6SiBSqOWGR4j5LXpP8rVWt3MXA3BsJ0ksSmlnTm3Aw0D0lFf0Ava2Y+sCHfIdDdUEOmNZn4X
5xXNjs//Wi4CobMC6dmi9B9H1emAM3cVzNFZbfEQ7+mJO9VV9VgCq8NsYeh91euR6Gnvr2qL5MjI
bk4v7p6N8Gvoq6/bgb8w6SrpR3K5kaL1R+ERvGz4DztYFDkj07NG7sf9unly6u1POoc+06UYCwt2
t+bUUb05CUH89+9vV0MGuuSZ9PnUpwK2Ty0NpIONd4je0MJhsAHfYldvfLeVbx7Uj6Wv2K+DiMxn
ZZxfR1fkKNJiRJRoYIz4urNh12qzHhGwQiGk2jS2lHqCNbCStEQU/9BWPDo8a27+/5UxxPVQ2EvS
k3Iy0SB3GjQYIYzbgb0kF4RZ2a2DYWp4ME4CDJElUoXlMtwsbP4vpPHB0BpmRLk5Jk+jULyTDNTf
LSV0KSrS8VR6w2KFGbFdmy+HNUO7UU0O4Iuzxx/3vCVDnGV1FF17O08EtI31OGeKAQBjxEWjPCFG
0ggnLewYWJYjFFZFgQ8k4oupDM0I+Lr7IHaeX1rOZPv61C84tKxT8TxgCB7UeWinlspH/ymypSVY
aKiBXAY2ZY8DmVKruz07c3/m28ig4Q+PPsjYNjBH//sZgFhx7urhy0BJlNvZT1WP3OkCK+ofmc+n
VSSHnp+TeXqtqsJqoQmNhjoXkTBv4hffflo/zSM7n/prElILmvmPstuB3Q1Q2SDFQnxjYPR1RQ31
gTv7lpdL8EtmGNArUvFtT0nvC78REldclIwP9MANyq7i+55zSpeVamRzjux65mGyp3XXfaqdW8vp
jUWFURQqiLXofapLLBVYpuSSohp9fCWcQMoGE86BFmcRM3AFTGJ1KFj+xfCkhkNVdBbBk76MtNgV
VXR2r1EwvC6Z1r6gVR5SiFbFEoqvcyay/Oi1dOUJauVNVaQSxr9AEfNujT6l8dJRblT0QIzf1hx3
72zjLstZALBbvRrnzB3pxZbBHET9FN/gx7SevcVRiINCcZf4lCDZNar+F6bIXj8WoUVPvAbn16YC
OAAIoXebfg65bcFyMh0qcgGt7zvmDQvzkqQKBCta73nUg3SBJXdMskzSQk2iIpuc+JGFvIsQgEdo
97bfbUlvanBBmpLdXCU9QsTnEwUKhq6iTbfkK4e46aFWDDr+7+GOvGwsuGbMjfG+W0IJALnbtOM9
iaMq5KHdgIclQnKX/b4lMvg4LKNxgFhdvrfWpb5JPfl+0QeRCBKjHgzw1ko6blSQZYqNG4mCj6qM
mxAPMBNudp5MNIKAYH6J21Ewit7lsQiZAr1MEMZDnXTx5Cw68LmcuT7joM2iFkWu9ak6Cqg798yd
MpzFpPhLbSqUJ7B/d2gNenjxKb8cYrCoY0TSd7KYSK8gmJaOE3wYSz2MyxALhheHJf4XJzpsjFkm
sri3dEjVVzqg5oCH8IHHUrpjS5tbVpwPGltssWyCpQ9inZlG/zwesaTC2B+Ea30RrC3y3s+tUzTv
HLPcx+43bOD5Ch8eYxXyIC2IX66nn8RK2+N+CUVz9/vOpvYOEv2O2pX8r86XxajR8dP9HKwqzxoM
osT7tdofdvE+cVIFmKYlI/mRAt2jdI7pyh/l5bok0gUO4zTeVuyrVYRb1GZniQa+kaNDp5LUWiql
J3QVkgG5pSkMhyEEMLfOnlEBn1+Gkjupi9VqWder4R/3woOugsF1mNQf5cNW/0JtZWMe2GMT34tp
AXv+T74od+jyEqrPNH3bx72CqF7LHKHQ2DjatzU3lZGege3+6rELVNMQvS7cHKsBLszxtUBJ+2Ys
pzGSFVpvuuIiu/VzNHqMGGvMZ4E8GL3E6qT+wf7bbpnmnpKPOJanQaF/6CPZMNv85G4hU4GojK0r
n3IxuCFk1CrmNrIMeFJ1a2hwXwBoa3A1AC0IGH2xf93dX0QGiPa2DZDq0FhLHwm34AexKYRzG9g/
4a2YbNHMJclo99cCdpIbXwBPZxOYUWzxhyYoBA92sRfljNjmtDH15d0RqCGbXYd5mCRbqLB0SylO
DF9xFXhr0XMIxUyVNAWzz2tOgGSCbkpSwrBr0UaXWEpMxwgI1huFWm/nlACaQflEVfAOD06NAlTx
ngWKY1kZef6dmf3p3r3fUXBRqtZEWGDfmhAKExIOhCEEZfSxC9em6yqR6YrjZhWR+ghpJ/z9yMx3
OS6yq55ZF00QhN16XuktWoN1fPi7JS/dsG39Y5BGf+BWWCZibX1xS7G0EVFg7YjFjSRUSSRTuETS
0D5LOat9oRiTEXu0o6u79AnlcKMlBcQlNZ+0YCVX5IwbFDQJlD4seeAvmcgLdY6957hAgAXAoBXd
f34CEGwA8MyNBReCjI3JL+mZRG6cgBqLvLSXW1NU1HbAYHFUIayq9RybsSBr6G1ObzN7wYviHx/G
Rc7HrBjabEb9SmnNb96ECEACSC3GwZE3zTXq6g316PiT/xWmt5301jYxbs2uCY/0WiT4wVEyTf4A
a2KPO73zjYJsSu/YfU6++UIEGldTw8T/Ljarsv3WyJ2m7WAeANnjH9whEeMtsqrjK8/WXnDkHl/f
sSTnAiy7rJBhB3trTV6thj2r0VIM65ZCuXpYth6ukwh3k5DKmSR4NVhw8PSyLFMrOSk7MlMYpsQW
Ulclnuf6F5TduaOATH37+HxIzn5Plg9SZgAbQIoW74VU3kn//CBCyePn6BLVp5QlvxriHOV/Yu7R
N+B8A8/UMDeCBG4mn2gtjJYX3ktcF+2JfabUiFRtEvPsj5F4m1ct2LUca5EgNZU0Dc5/3u3NnaY0
tlwIAWM2/oGcCYaJniEzpBfmK3CiLU/Le+hojj8a3pmoJC0AqTNpHo2AQEDBOVifd8JDlrAveH6K
BB9NGLx4sh+gcaPb/MfxrKh2jF+j4MY3QRrHEb3J59NxToYrRCvJ66WemtxcP4P80mQkNxZxRgH6
9CcA7+5rk52dIPqD4lC4zW7vJpCXh3w/2wXSgVTzqxwixJaHX14FMIBGoURSMHgc8r/Tffnb/UEA
mZw2geaqBHH6S3OKi8+0mSTl4Nuf50jHRCgGDk5iFJfElZB7l8KhMcggXaMmJ+rWrHIyR4JrWCQ8
s9hB78Ejp1qD9hpOgXmyoDdJHx8eFXYxd6JmZBEpnz9/y9o2YLhVOTw+QuaGYXy37ObildIeMvR2
4SkSx7gnvffK9l4UPquurN2ERuXgcpxQkhlIhukAQlUJgGjTqnI3wAtVzfZAH+SJr7uFtDAUYUS3
DXwM/UM+muub2yNpbAkxFW6dUb6vFVXB8dJPq2mzUsU6hMVQqwyQ1YknsDufN/FuwrsmXYQfM7JE
so1mkPYiy9DFPVIY/NkEMOxJ3XpAphjuK3Q9+cPUQVC0BeEr1lRjQpElnJ0t+dPiMzjyF7smJdZu
cgtB6ASxYG8VJ36nhd3zfU7cyRpcZSVV7TfzXwfLsyA8H/uH8o/hRkx1KCxyRDbtlWu2PzwFLFGN
C7sVV6ERBPrPoxsPnHZQwY5pg+nmdltCBPyEoroHqGz7pQ+h7ExuiGVUAxyn2Nz1dHrpmEogH5JQ
Wl3j6LJNheAC36x0VkzXs6D+paHYVdRX6dJTGVKslQ3j6wqp2woC3zJ4DjBh3YBwGTG9X+WtAiZ4
e7KZ/61Yx19U8xSUoTSnA5xZ7SoVucp+Oert0a7mJu9Sr3wvPzuK1gqhA8UgDH5U/T9unh6QE3g0
GslvbOqLYHNlNjhK3AtPswFy+1Rejfguex+3yilN0OUatfmcZNy4UcJ48t59qH4iBLXlF+WYZvvD
rXVi3V0F1NEL80OazjF30/zFHpmIPGhF1SgKOpu5CxQpeB6QJiO3umIjL6tz+f9qjNtkxX1rs0MW
aBPCdFJVBRzjn7TzLD7VL0bqoDNoA1pmFbK/arlPTKb0jvygMh+vb88llk+fotugnylO5QEt4x6f
3+8tnVxfupS3GkpI4mHOS19dzVeowlFBe+jSSMNI/8lRAFOWblb8fbARDpxVf8rAEEFfABMODuKn
j05C5f5Y2YdcP6nqOEqstmk6wldByN8Xw8YMu2EEH/YJkuk6vJJLqUya7O3hluqLMS2KuZDkIueF
osDSXqIjxLHIWZXXadysXQW7qOAA4Un+LQozcUv57oahuJ9NFcY23NcZ2ae3MHnrV/fjiveg31El
1BmBSG+EqbZPWjKFcFgReKsVkit6A8TBVTNFM4vBfQV+mfYpH6+nOm2XAx/gtTx0CKDCFMxdVN0e
XhGUOzxyY1YQDZQy39kdMYKrLBZC8PpoaudfCIM+8r4GXh7nwKt7AbxIKSx3n54xTeEq04H6w+vG
KP55KM5TMpiYRzsvZWZQWN4Kel0tl3XttftpjZ/6qM5C5bIHpEpuj41do0322mxefpxYwpZKcOrG
iPRa4ZtBNm7uXyLEm9+2rtXXRQuvWQQE3S9xeDyeSXSgud04LXnVTbjtekixZfwypixgMFfSc713
9dINUT61+QwpXLbnLTWo2zMkofkNPKXB5/Rf9WDDjVVPRwDBAgXYITcCeQzcAQuToq2kauIHJkDR
6BERRZuDSGRAUULX/PqAgijk1Bx2UEZ5qyd4xZ5rvgeN9NxokOon568k7fHB4J8n6B8VHQ4wOsbH
a0xgfycLHvzs3XkSqj7GjeBcvwJivj4m2IfFQxaOtkFEiLeUMhcYPYXcbiKKtdzTi96JLF9vjRV5
RxQvtmjknsS08k0IPaYHPhjcbZUipGbLQK0wtUPGfC+/+jPfHYpNbyXFcMTyaEyA6Fw3WSPIaPWm
rUu6+xit7QaKW0EYE//GzTd9yOb96EaD6SeLoO6OmYre60cfX4Nchrn/2iBRIsERLy7I8W0crCz8
WSqNSqxt3EoeXN0VwG2wytl0H5XIlJC0iWBhX1cIhkoO53Kz+Tu6PU9wmkRffnS8CG4dYZduiMbd
+zWNocuKdf97ul8mygCH2dXp+TcNjCWXs0OFdF/MUiU68/CZGEXAh+3x/KuYjVyaejVGpnWEBF6f
A2UFRALUmLltqgCNDVeIjycdCbZ7UXvhARbRxt57StnOFBSSeEAZy+3musrAhxeTlKQ3bkCiMW0t
cfCALuphHbpfTyKPGwxstNhULxxAVkM2HS/vnWZuDcqDQ+047SBZwKuy22brfyk4ZdP8lKUhsn4t
uKB8bfuIxTHH1cJBe1rJ0uIKimKPX2jTKP2EPoGIOxS+PG068zWTQe4BAvSxapI8DwYzHgGCznk4
9irTnAZfdtjw3xqTE+qh0w03fnUx99cOOxl6ypsvcfYYZfY/hCtK+GsZ/d56FTpj0czUs7E6fTqY
buzxUPwTCI7QmbIngnR+f4RvH9TVjtzwnLZj7VmZ1+ZCFZdE+D6wOL5hR3XtvSCRT4jOY3L/SlO8
5Yd6Pq/sm3aRANeYQJ60sPS4r0Z8xH++ZK5bWE1+1IPry+yvn8n5Xz/PDBH24j51cTpw0cskeFi/
HlR0H2ls0ahFmyv15YO/ZTXFZav0fV9sN3Y7+3dTSX+g4MT5NpuzKZYYg160hkOP9pEqYX7MZZvl
J4dqV2oOpb797CvWOc1tqWzpT5pC3uJQIkFkKH2gf/3gQVwO5npanf0Cqz/luyXQmRMJ03uXrMHB
CvHn/Wykg/DQqxsauJW6CaQYOX22BITKwsikst3PZjWQh5HEdRbBlLEaVRWTJSCufZcGCYAMGCgR
jta82eO6W20tMnkr56HQUzTv4UCkbUQPEKTPlV5VDP08aotsXGPrTME8gtTiM/qAKXZeQsGoWo6Y
opFGjGBrhDr7KqPyGpF4IHepjVUQad0ujxUU3H8xd4EWGeguKqDMIWNtJHRX0oIUjtXJ9Qs29xY1
olYqFrvAAOM5hMtGyHo4UPlUFWWxYOuT73DywzM10oRTUKB1X2ipppQ3NXcqZE+mZlOU3EjVlrJo
2Ix1lCTnnmKkw3/IGLxVQ0mehSPR66guPkQ9cAqclGodMbKznTI4nmjpHz5JdEaCwxFvrB0lcAgH
id7H+lnpZI2I8sjHFlmb7+L+aT/4lZG8e7/uKBExDvoPmrwm+U672CYw1TcMOBLC63jWLLaFpb0N
j8eVnJPJCa3io70x0+cVfN/EahSbgvAZMoAEsuCNYk4kCJj7TcmbP1/Xx6yT58Y3ag5urUCxFJrf
a/PGG5gLW1gx9ajIHSo2dbFl7EXdJmJ7iGeZS2Loz/5mpHvWZb/vBJ4mMAqLggIMw2i61n8OEfVq
184lOu5gX8cuu/PTZTzBmtWfhPpZj7lvI5zrt0iC+PugH5qBcb5kZE7C7JzQ1uIHyg7Wx0SkfNGP
ycr8tbCgLAoy5xvv7BtIAZQwxsG3gM5u7R53Js2L71DJor9LpiZBErnD6jm4TlgUWI7itXz8bWBi
OfhCSwCtbDJnodqDcPwDfF9gaZ2ZzntlxRCDqfpzgTGu8lBdkH5hgchcbRzwgDsJJg063kKVGgAU
ie17mgJ+ejn6NZ71mJMNsIWp14r+UXMk5wOy8eV30S4LyneDP/RJuk0NKygBvWM5lbqkd3VcJixN
Ebfe2lLsjvS3c1sHNpAWJ73GRFXUQUKVfy8pLdVVdrvHqUw7Ir8mLf9bBSq1lXTIRvOiULX0YzeG
tEm7asXkd+u6nYaFcl16Uq0hjBpuH+15G54eBgkaY9LYMzpL/qdjt1HY9Dscre4pE2j4fRsFIgZz
1y+IjjPjXqL56arAzE0sZvzOFNLKCKu0k5hprkwgW2D+Bsr4uuBygPpTXku40oHDZidPDn116aAk
Q13kD5+ND8VxQbEPUWSVAS76WdPfx25+b1OLCBVZRBdIYcbCU/0FBC9BkMNHZjaM5vaYlSqNNSMC
AMDSI+TbRlls73xwZmuVuOnrIcTJYhY9+f29yeuG2OcPtJBMpWz1qyCUBxNcrx7uUc+AdIBekRXy
E+LrDkhTPA64Rzspq7b+TgbcoZpcNauP+qJxhyLZFMOSlECuXMuBCyh2TkYU2wXYzNDKXkZaAVGB
85OBJ1XvGdzDRsrm+R/ByGkMS9HtOIiSpbmE4LQ6WPiaolBvSmBz31AYGfBWefdFSlAy2KT57Gcw
9YUh5eLZ48KsQD48G8uWH2gtUzLBGydLZIVD7X85MUSbAReSUfjg4vqeh6vHbPcWCBqY+rYxBNye
TmbO/Vp2vPYrKj7I0Sus7PrE10sQdEUzDI9FjQqK/N7xWa1PQV1WCPXDzHKn5b6JWoFu9gvUK+jT
IeldhdXyLWSvIb4ixAgoDaJpIKD26ZChVl1cNO2BJhp8c2bbtFM5ujNKfmHlBdG9WvGww4cMUyzk
vnPRjKFOJ9pQWaTqHets3MdWHBKaR+yhrAfYbbqiWQAyf5htkVIeCFq6flVNaL8hqI0VLMVKSoSO
XBCjmt4bDWYPfkxtXpFTVyiPjDj0U4X0rovrWb0Rtk2jNUHRw2Jy6smcu2H+bexbID/uTDQJETmQ
xVVbxkthSs3LzjmE1vjD52uLEP6ueERlX5DoHYu/u18z0rBrqDrcJlyUtcDP6j5aqVTZRdTk+Ivv
ChNZBed2KgcVt8J9U5XWDM5phYuFTGR+Qy/MAU2L+AhPtyddobjWQgBMS3LxaJyLQpiG8d1WrqP0
fNjaH1F7A9VmZuy6tWDVj7cynKU/rWiLoDT96iGTiBfTT0JVH/r4dfHaLZ+HrQ6Hs2m8WPsdM07d
tFb5RgDJG1pK5OBM056Vy/CeGP7p4E0Uti237J/PjzKK1tlJbiT2BNWf0bVH4dIYQwAE0osySMxg
0gyBQlaCLBgP/xULNHFdJ7+s6pAaTMYlaj4maFY3ZhIhDvWIHd4ZYX3MiliwUJ2H9nsa9jIm8MMO
HLhmw7oeMuhMvdD8wICI3gsTHbI1S0AKIH8HmqggLaEsSYroDwqxJgm+fWW9ykCM5i0A8NFEKCAl
dLQRScB4orCK7uMhPSfTTLetA5uF7raUXcvXoggpHQvI6P68oIJDnZrNCwwdZY4q0OP+fK8Ngss7
SvalZqCinJD6zicupB9AL8D2n4vM0aEYcH14BhCuGQWZqM0ZF0bMPFAseIJnmStvhYgNYGLjUo12
Ln7lMHwVJQNtafiP22W//hPTwd0iA2MSrXdM8hpw8LTQRmwwjAAlMtJ9iwXj8g+df1SCNzm9qxAU
by31dXk81KTlGmVJnLwPBe2KkjVbM7ext7M0qtaebsVU6+vz3wRhDdAosHQxLGeF5WJ7ouNUJnVD
CM/za38Stuaqhg13hS2WnS2yA7ND01+toZqF3F2G23NxlIvc4m0t9qCf9Ksls7sILg3A300Y25HA
RtqC6St8qBm7OC2BWT8kOHFf7FiZU93DGWARf+rQnixTqExlyzVTret6DKWNY8cOeMDR5sULKdP0
7bNV6ETUYbvWlyp7hIsagqglW75w/TzPtLD0FBBVLk9iSLJ1H5Lomybu/OOskJniR1mt1yx9xjxT
Ev0nf8LNaOFRpa9+FbtWrgXa1tUz+aDGpRwBcbmN6l7KrUZPLcZhfQTfUTiowMro9CRqrXKu67UZ
jcMVRX21kI6XwVrnQZpWj3F6UNahdHxDtZggB4P1U/YUs4kOtP463x9F9tVqFC2gmVxUbZJW+NFT
y+U1swLnfj9owvkBS9qnBrR/ms4y96q3Dc1QZ0VdmDjBZh1j8VQIFOaa9U7Jk3rRBmAsO0+pV+yQ
2d4zElAHwe9wJUZBpV6rJb3Vwan3Pnt5LOw5kqoA0c34BsFbMda+zPzt2TWlRvQ6FsiFsy3dE3ET
vso4m0X4UMPC6e1waTKFHURqSN7ZQ4hCqLLVaRt92MONJ6ZCf61VdtQDKUFyQaxlq2wTqOgXOD7z
BCEQRyV+c+0e+aP6RNPMRE4LbCG/tErPMwm8g0IBDe+mXZAPR0D2uIQ5MWYRQ0dmXlQnsU11cmMB
lqn5l7RRvOKT9z7JPvo/2cLQWoZaSsj76N/zT3a6p+7O8SOtTGIIEBXZyftMT3vc5ZcqssI3rGmA
dd90IQxAJYwWg/zBas+TiWtwigjNMEjglgIGG6D5nu0kEfxPWWZJ3K5j9uV/eoTORl+4k3w/F0pr
0S0KTepUmzU/AMN+WjZsyoRF2Payhfo0W0Altck1Oc0uRHU0NPBiI+rgHYITm6iYUDgKAclVg7+c
h1kog9Fq2YgM2PHCP4nlEf3VGrnQq3LaFrba2Q1gjbunEAB/ENlTiIHoOSQ19vdOEDvoOAf5AV8V
bUiDjPixEGzOBN4yo3wl3EVgrcOkPdRH5/9UxCSfeIh5AZTyl5XtByoybX3dZdem/yr/CbUXimKa
uX/wAQnyulDXV1v5k51LzlTAFaK3fomDWdyHZlDXBAYHsZpQNW2EFZT7KJYpiHN/brBEomcNx7pU
6Vj74oag2qPox0jhy4yYP3+qngIXnt7ADJIU4gBiEX151hAx1zsdkVUMnO+3DEc11RfoveaJx5iO
D7tQp06zHO8xYynrj9klKW+r5Z3h1lP2hm19neJFX2PuGY42QTKQ+QsDQzlSD+HU/guW8W9ZbYmZ
PbgmGVORSDZcYzWPnO/nJezxGOcB+gCZr9Nn+sqx2zri69X11VYVtFGccQEwfnm59kDUV9ser4tU
UgxvguwafkxaweR64RXfAoIoC1QsE409/qSHWMiWJkKz/DmDAnK0/4tNRqb0EKnApCgktXlLGHNz
pN2C1ACoiiprCF58W8Juath/KHeXsutRmOk7Zq7rx3b9tAeIfvPcmuyReILEOjgA1UdFhG4leqjz
E+dE7jmD15FtXKBkApZNzBtu1PHwdUhVhusyHf1zajJDiICot3un3jbGgJlkuSCw7EhGGOJ7kQuQ
cAv6NyFwB2VN48fkILZWGq8v7pCcVOGhtA8oBS+LQ2+MUlT1iV1FkA9ZXBK74y27In6UtbqHf/sr
HE+8djW3v3av6Lt2/ikthm29ye/KRlZPpWtI/SDSEQMoQMmDVpw+z/COZt/XQWtCl4s1c0pFDPm4
AzdqHj/zCTpzPFVjq5jBJyCI+kIULqD7oZTjM1ubL2b5sczz/o8cyeBM5olmjx9JjQHOTzHCuRDm
DW6xIS9FVFTL5yCCYFx0hqGirXxuPFpytPX+vlwAARYOGcg+68EchUEQIFJyl/m7C4kcXRoz6Y6T
vgbE0601CLrAkbET5UoeGhRAnHOzvmllYizYE9EPQoXpSdpzzcI6P+BRa/BX1t3WNUZzNlusZMFK
aYU9CMT+V7uDACzFZ6yb0Gd8sGo7DYYnck0Kp1iwRVcDRA3B6Xy5ZSrwQgmUslQi6T6ELYSdknlJ
66EKD7F3xiV+Cc1rdUYp9mHZjNa7ufYWdGF7xnAdvKpOunj6pWRHBkQdpby/qx+4gcOwMhjezTMB
vdc+VHFSpOG4674ZxZHUagSXMoHXInRIKFcsY0KJciKjMPZfpgyynPbdSbC05PCZMbMNy4SRZwIF
mUEapkadkXtEY8RmhvGqFyIJwybLLdOaCuT6J6jIPev54YVzF1cHKZQ7G45a4DmiiuKyw8Oiw+ZX
fzzDAoLArNYMFP/sIk4iXnThBkubRVgxB09eqlCnJFLV5xRWrSZLLC63QjgKK3KYq1SQ8lyh/dC+
Z61Rhxvds2YZ0D1WL6dGthFz+35DHDhwzgegfrtKLc5Wg7xnaX4xXpmFQ/ChHndd9MqN4F3Sl5Dx
dsyP+QNNGM2lmWIQCOwhQ8RAZrvepvnR8ZY65flqaa1ZZ1DSAwXLPiZNJM9FB3gu0RpUN77bOYBs
iqmaQSvjQk7+iX1AwBQkr4O0FZFXmud9JutBCLqCNcpaaa9ipWzBMoeCwzf2Dug7zafBVvd8kW8T
cTvN4dXjqbxnlgqDCU/Arvcroc/1sfryA2F8b4jLZ+a7PNk0b7TowqV+6qGGax1q9DHMIhIzwtQc
HPZvM7JVa3a4olJ8HRcUrhnCrGFZ0gFE/E6oXba8a4jHfVkH1CC/ib5yiS2FJb8fJXJO1lcanwp4
e0jPJ3S5jQnamudX8txSUNkn3mDMrdvEWJiyN1mtNUR9PtKObtEeksS+MPWzMpkaqHE5dIzLJnrD
sUkbwuASFvIJoj/D8TqK9S9NYyQhGVVPmlNSP66Ut9ys0HhsHObOXiL/hkoYFvmsbWwES1blkFyT
OqnCpvEvkutJMDUV0uUb93B/kmlVGP+essKlH7wkD/bDH3ttE/XZnTZxREl2xXENyEgxPFwo6Cab
Rfnd64K9JaO8RerLVq7rkOwNgBk+vxlsjcyEq33hczvl0mOC2fE9p58l77uZ1tK6TJRDIfKvqS1Q
Rmk/CrdjEhz7hFx7mVjYYPI6fdQX0xzssOJVmh/fUriUtb7rb/FKzxgBwUmoiMYvitCRQdW65YnN
6yfKsN07cik8CeULW6zVgA0B9oFIAzX6yPOijh6IrQzKH0+FqVoEaYXsVUwvmRxgRv47fXA/NYT1
9kju/NedH0pk5aj8AUUr1FX4XSJ4L/OVWgSJZouIaDhj3Vh3ISno7zBozRom+770MpkE/ves7TcX
Ovk3sgKbgnHgfeX/TzlPL6SUyMjI7GGc+QjS+2ObCPqnWQrVMcJpUngXJekRobs1U4G5UE8hfIeo
8UDNUDrXQuQ1M5j6wFEkgwF8Z+BO22uzSKUhEZOhpE2wWZZeB34gs4Jhq2gIYWslR582EMwP1blH
RijTtVtdZ2hgPrwPitz0QUYwDu140AkblhliGyNmdvERAvqizO5E5YmyPZB+Tfw0kPr31i2oEbAd
CEktVphpQ3vpqrGSLgl3L3MP9txRpQbIITEfCFL/tCiwp3sEKjP+IRVtdqu6UrUNYWkta2DgGa7U
OgxPZ73FmSAntswnCg4wQE83ZStxI3Lr6/i7j/Hfk9vPxnpuTYO8qui/0/x9q5u9Q9UjL69o6I3x
zSB8l3dT+ssfkVUp+8lDeX0vwwWl57NZNNdSkNSG6A4X836zRQMdxDtA4P/1i5JY0GYPVEN/L6mf
yfKfFElZe4IGY+VY9BsZyGFZtRB2SVp5cwIPVxcXJiaO9MFdBiNsgJonZY3hNL3EMmUcdKx48z0r
JfSpX6dWBpLUmfUX5SjlHfNCArbC48FGXMH4A74xMDH/zK7F83GMqnZcGWRihsL1Tpuwo1dDSztP
Nak1azzIVn/QM9oxRjDa25VQ77AguX8Fp11gNhzaLz6PSHlxbgk4mHXgmTiEP8GIcClRrIsXcdJX
oYL6tc6ZqZ6De/gfpxP3WjvkwiLja+Y0jXokx/hEA181tDlNIVp9iM263v1iuZ5WNdSCYA1mO/P+
hJHjABT8INinX6OhAya392fvn4EokXH61VPrs+4qpArrmoOqyBCHqbaS1uT7YoTHZqZCH7fGCouR
+JDnWmoQS+hba4gH0Aqny3Cf6V8OShv29CkQmdwefoz9ZIm7yEL0lILF5Qq/5gTBNqFxY4O54mBw
PD8byHL0tzBzGXC2viLjeGwqTJiV1VO8Wr4ojZHysMlW0PEWczgsLnGg8X59j60y8Ib8r3wwVKBf
Uc1qihhG9ni0m5BjArGzNGOZFeFrazq+uwEGpvhbLylAf72V5/ITrgANGKpHCMbsXTeWdPvYpM+3
DfVUJBj3rmfLV0BDvJIVwzdyZiPvK7cUO6B3wyHWWTlXKvjH9b26SkmrQa/iMKmqoHQvMno6/Emi
p6YD05qVh8Fi704fk5nC5aK8P0L2xor7s2XrDR5au2Ob7lviRJuQcX36LTpyN1sq63MLaQehOrio
sY8EDPl9pmQx7blWkkzlRXVb/h12wkHFZQ1HpT0UNVDOUm+4DFIkS7QuV/EGEp4KiYClAukfJVs/
OMTREG+dLfe2IoBxqthvZzSmfSVAYUPEbFgLX26B2EEHb24v8w9vhoWIwcvUhVOsHJFqoLhdm1Ls
hyxu8xwRW8N2ioWNGGzGPqFsTRPx0p1lAnJlt11sWVKh/FhhZY/DRjmHGRp6Co97cbnpl598pFvv
zYHyoSZlGnFMoT6unAhaaZyVoSgiuYffwbV4R9NyIvym9ezTXcYdHkeURC8tkEy/q7WUTeL//79L
lbCk8dLQY9lmUqgo1lVPowmccMYFVzooJLVC8hRm6egPxUraF4UCAfdoWFD8A8SKxq4tpigaxZ6V
1XaCRHqSz828pxhuW5icPEAsiuxa3gG1hre/DvphaUr1z9wFsv/njYwFtvIqJXZ87z9M9aep+Hvx
6A5BWi/jQO9m3P+DEoN5pCW0R1QrFBfuH+WZsscFVPIM/KhZbs0gV/P434tavMfIXT5wKasnRbWf
hX1uKisWwFjF/NLbSE1xAbHvcUDLCzHgSQUY1WzkpteRnVQsV3uauBG9/quzaOi9xMx3ZgNUJPY6
da3qRlcAiEF4ayZJQy+NML4vkEGaMD+MHUaOV9Q5Co2ODbLl187+PStcd3uj2A+0j0KMPlv7VtlJ
kbJMFMDt9ZHBAgeno8uwGIJm5o2OrBV06au0Uef+AKs3MJUEC/84e3dNOaZDOqPECqPiz1anLlV4
eqqCOPyBL1dJWCpWN2xISbkertQRHeBeTYODRmjD3hq5dHs/UKDYvZ+o7kCkx+mf7IhEd2BaKsxd
U5KgmKOe8yx2BIjB6ghtjtynW21Y83ix5cnWz8Xxi2UWMOStwZ2hnCoDezP0s2aB3f2vVRumbUkv
q5It7V1XTrMO5HF+u+c523eM5quG++4nqrXT9FtnSq3fMoG6Ml0FtlNCEF678SktuzgAmsZZS7YE
v1UR6i7teMK4IjmZKGYLZdSQtsS1yj5R4DiJVXRSKRoZElWMBAt9R5rOoxU9CRPgVUmUCxKKvlNN
4CsKUtafQbyxgyJR70AnwY84agUKq5zJKWtxnG216dYfZeN0kEvuGXgna3oQE4Gw/i5lmkyAl+zm
NFpDUidCfug738obtR2U/REfgl+rD5uMmVlCJq1x83SULWBQ62L/rmSOoHHrF81vlDE+yzjDs03k
vGFSR8t2QIozHLLOJcRjhJoglJAAdDza+b1hU5alPLc43g4bx9l4Bff6LHzp83wq4tm2FKhadw0t
CvQsg3zRmqiuLR+SbBDNP76xg7ppE7GC/Ifwig9csPwFnW2nwWBw15rRUJ2TzSbR4uTKhz/UOh4D
drhVICkwRXnGJo3NukJJ4EiE9iJPdHOy9lbZwz5WjXU65H0kJFe2MEFuk5dZ4oZ8MbYoMz9e+sr9
0vSGe5Uiwaeaw0e2AZOzPO2lOf7+GA1szYI1mtQlswCVYtkOubDO61AS44L1VE8TWjthzE5vubUS
yBGoNih0NAM74ysmjwWJcWDf/zSHfzz6qX0EUsvdX62lUitbWf9Dkrhv/OStoJiVmbbuv8u8C1+K
4XsPoAt5Y1ecHSLwWzviI/KEtFlCdbXDIhUOF/pTM13k6SIrXqaVJo+RKjRxdaWOkJn/lDUzJ87f
bJ8IPa8R0E6uoOXQpVVdcJxpdekFC/ZXBTUrlNqYgYXEUAEfTLBZSBUkMsaLxiue196XsMG1gxU1
SHl41SC6LBQvyCHhnqHGRirYIaDQnfGR4mDYt4YT/zNyLxBNQAKxGmPEqXuuFo0d/4hgs3OtWoAM
0GJjPO2uf5w4SNb+w1t198AskFklJkl74osPcHFv/DhWehymeeNNr7Hxm0JeyGZzknRRV5yBG+n0
pOoCj02La0h3DttWkEiGudrG2HRRmt+X9HzMRhhTOiMnSeGBwGz1Q69ZpmdqtKiTarKD9LA/4sp6
gtRwGGdzLlfH93BqBBl1C1DS+QnYoIFykc3Gf1185uXXEjxENGbfxw88F2ACpREa/OCa2Qz30js1
i2ebh6hDs/Lia9q/W4WnJPyhAjGGr1no5va/2Nqjbjrp7p3WcTEI3jQHQcUwI4zqkOT9eUP6iMa9
MzqnDkCFaJUHHGNwl0LMbDU4JIprKw94F7QHgheAxBFZurPhjJM1WjUBy4wi+G/d6WaAnUPxqELs
ZhnaUEQrfq9rhAuTI/MDVjgmlhk1IR4pskLdOlCtPi//TVYA3l1JAdbjZvC3FY5hrI+FdF9sgrpZ
ny7Z6C10aTbyLsTkHFzFdB7lOEfGeBpJ5ZxVmYTwr1oAptgyDefYcVjJ5VIeHU2JsXBSI5tQvV1s
JF+FmHwGYZJd2Ha4TDjmF/sCcf6SUd+O+Ekfx+mZfu7D93cniUw2Dw583gYWpnAajTW7eYQKNJY8
JD0ML67qjrmQOEVHU8WcgMhLm5M2xFW49HKsr9PsVkjJTAUUkXoVEWVR2p9MHSHlSEh0H2fZJ76O
9xYgBTMVPdyWBUUQRLVUyY+JdsAuCWoNjfzMI1hJILPlhbxHj7JkSfn/ZgqCOlIffPG7YucrksrN
oXsK3Ik9YUsHFGH4TrPmIxTtE88CRNKa6d/UsP7wb8uwtcAoSUFN5dpOXtetSiLkn2eoJ3CSE+5D
FOUAsldH77+lYmjSaPhG2Mz2svnE1QBHJl9/AXx+gjH0Zz2RJNRz2SXEJOAFeU3J3YYGKsrqLTrP
V1/n7fMQAyW5czjFu2j9/Fg6m7XPyXRJ1NhV0VRsAtivQLv5Icl8l5stXGkaZaQHY2HYgufrVMgK
wqh3pRHhEA1k9Zoh0mjHk3n9rkecezRQozJ3anxxS6uXxCGJnZ9w/wmDuGaqHIY2LP3gdmxhp93c
EIrvevoKH7Q/+iykxJk4dr7FWupLY0QrwJcqZVHdiriJqqDu3Jvb+3z02eFtKM2wV5OFx87w8pTE
deEjvjn3HvwX5PDnwx9vsW+9LkvYZ2DfmUodoHiQi9qO2Rf2iVlRY+agvGWTTRUvjpVCKci9/51i
ajupXXOCms13nrBpOk2q2JAQZT3vp7ZT2iMz8ZEvJY039CsMnDhssTZvWkZjPglU51ugcIO/dnaA
bUm7elF2ocHAz2L5LJk7RYyybRYM4i0lajI1lQg5gsZ/splvgOyxh67fSMPoUFw60mEP+U6N+gAi
unT72TABM+g6AANkJ7K4HRvp9LT/ic/uH2EuuNnu6IB1ff4cA8QxiTQAw+a2/j/mfKgFtgxIa4lg
JoJFZTw5Rd0KTLr+N0oTjZoWMoD+WnfCeZcToAN7Ath5jYCy2kP+PH/hnDo4JLCWMrb+OaXAa9F2
HBfbBDRXscpF9DSjQqR4YLgg7KkRzz9aWCjFSNoB0VmB6b9UiD2clwvq3lB7Orzv8v8o5lTv/dOE
41GrdQ6ITHClBbQEphA1xDUKpIB+bgBEAfRGERC9oLZsLMZnxSQxim65HJMvCPbUsGEBAA9HuIJB
UEvUp0rB9m65++KaN3dmEsWCzOhdzV8e1244oTjiSSHnXzKxoGFItiPOHT6fkgiixg/AAssWOCqp
oJufjcTtd91qYWJYnwvAewlmfgqiTaJJgH8kHfpOe4SViYa9zzeu/dxgZepEDzD2BJ8G6wCuNg7q
v8QgzzhKY+VM+bMd/tmA9NlNtVRFVBC4xBOBxK3GMbXkjLVOgAz9OulJvRZg+1Zqon5Ts5Y2TJyE
Ljzyks8UVkm18vRSiMAKd1FZ0B6AQLpcnU7K/Jkw/cRNkxdZjx4E9x8jKRo8x3JjO6WWMryYqZBX
dFPcf4T36VtW+K8DHoawNUNTs4vLwIQmi65z0u7A81d2mFT7i+eXec5eLkdnnD9Uky5wCgwQoTiC
4tdYlgzXaUZR+eD8Nbxr8dBoOka9wNJ6y6lgYrJ16gzAj14mkgTYxA3CGk7dD5hTNsHy4G5C+G3v
MjX6HUjo0fp68Turw5nXlvEwdY7Rw1G47HUkxJ5bfKiNIb8LZO/EBaD8EzyQEaeVWHbGbmAIogej
W3EojXmSnEu43kghTj2559DTazjRhVuAeV6bo58+jVopqLfbh7wk8YlXbG86dDzMdytdJqTW1SjD
BVSwyiEsu0DZJPzh1YBW61LxXGZ9/zhmPuAI4JfPAlOiEmeBoNR8fCkIEJKgWS+GWm4jcC6eAWfC
GumnK5aYlaY7m1pSH1vFrRX+t/+dwvVzHhSu74K+27BS6LISm8tUKY+IgkoMW4dem4skWxOSf7l7
eh/0sJ7fRzCP/gU81UufQmTfbnFytvfiLSHN7wo53cPwS6vzU8D+7WIChMhLRORHCDKTy3Gpw9hh
mEXfTWtkMAwsC05IzjunIhOYTs0irG1yVL+coGB77dtN7ozxfKUFf2HMiXmgTA4kXYAglt+3g786
lX62W+8hY5s0R13MBYfBcQkQTrgcwHVpjfXDcXuPktC/c1Hjp2Uq/OrShFYjhLYVgJq6YTr0ixDf
nuV2ebUPfxt8V06kBDKkitFd+0r8Va04Xl0bwSwOPvq2I9EkNSvhnTupi8QHJzY0KT21JUu0I0+o
pJ7F9Yntd1OInEI4fx/bwpPK2SzfBqYH0cyHlGx800IXz4Fiv5Usjrmt5CBAwhDgXKaMPXVKLNVu
6JaAO3Rp1wSIEgfS1IQNe4e3Pl57x3uJjC5AXIJnl5eda01ok/xIALvseZkG5BWmE2eas68/m2Ez
KKeaAXoLEi406k8KOp84FGudzpnv9O9MKD6XM8Url8sa9kKG9mXnxPlQE5zW0st71k33wnvInF3P
oHJ79bQCJxXhSY8Mmy/UBdtwH0dOrYaKB4hC7t7Zm+H9juDxHOa060h/uRRc+BXcTL6TlJe52fei
D7UezV3Yf+AsK6k+pgn3iHk+1e4rDboUaIKx1+K69WPb7+cS/YBNNW8MmSvkfX1Ps8KuHbif3dhJ
RMxE7whYD/HgMCS7rlJqgtjlPRYF5PCzY9Cva7vQprdsMInws2CCTFp5XmILFs/cVURkH25w/sP5
JjeGJol1Jwv12edkj8kr8fVmnxc2QBRbkPw8c7+s9gMsZT0jUFx3vnds0nTwhgCb3+JsZnpQnyfr
ijWsaUtPfXJKDVy4LvBW5qfQIdGk2is1zbXWtONn/j/siMpDJPWg19doJ3YRPRYfYIGxUKsRUCSq
pBmuJ27+Gw8XCvm/A/m1wz/j6KSUx48ov6p6bFDzuuvW0Aw5SBew7Z3Kkk4/tW+Ef9kN6aaAxPxq
i2NSTWwsfMRM49UR60FQZ3dInXKLxSjUirNgpfRcNzi5VCSEpJtDjFsVf2MfweYP8655PqvTqqUs
CRVoUxmitnhPIPOyVKYbX62Y55lkz1lPk1RS8MkZBB8JtmE9qeLUSjtnuEJAMZ3xAj3ICERlJ+I5
im3HxtBdI5u8i+WuN8iDGgXVW99FSRbcwrWX1eH9HsujvHuDUCUeDABYIWD3KDJ0dEbvGpco+1V2
0VCuBjgAx/ShI1DIVJgHL45X1PmrRkk2WHYC294SlVGAx6iT/4t0hPUZNUJw4VjsySM3gmfXcm6y
g9sggcZ7co81kbdbpFkuGQfyXsrLrNEyjL9Zvs4iIzuvwpO77dKmRuoF1lJGkGhXNntSfmBmT9Rl
NXN9xMB7tTZ1q7jX7zNvtINWlRfbO5HPmAj/PChgg64B1PDTarYaacIDA0UsWVNBBV6eZhhUbl1v
NulYqZQxfA4HdnbLTMl+WSW235G8yDB/XWI+U7Or2snvTOKJR8tqNJbBMk4pljMQ3YuEQe9DI2Tj
o6KUDBsklT/tg9M3TvhfyT+6GDj5pYT8uE9PPVwddyuuy1esQ6ccSwhIUl4AMUuRUsyhPFkzSnX1
XNlVmq0g8MKyEBcI1wabQ8ZHjD69aS/MQvpvPFavpCIuYI9H1YnEdjMOUcdwL9cRgZ+vwrOLGWOP
NCyqeLmSLrye/0jWSlmfzSO/ni35XYTQl/mDUGNsyMAbfuAjcGDPJLkmFMgz0tJspFsA8exwXEPI
T7KYmo4AqE1//rkEgj0zJ4Qhv3VRRqdIt298LEZMcqTJGX1O5CoTESNCmFtYGOA1RAqJ3G5d3knL
5RvdZbJOUC2ZESzrPoaLuVoI7kn3q1SJkkNCYrrZwkDy5xYMUr6k5i1E794qQWtmt183K0x9nejy
JomNUWHjwIBqu5mBfoaZ8BL0/SpQVO4ckZttHDiDYmlijRDSV18bm4Xfcf5csuuIxApIILOg7h1S
CWDdrUNyb82a3hkcLW+bAerUfbHb+4mjnsu2EDhr96tSeG4sLI8ygNGiJdLB3TX/mtzTtpSWjKgC
gFf0Dp9pDLbjtNxFJ0mR9EEoLj0aUEvVoPXb+QupRl5kh0LaqkO2XqYGnSTXq5Jk9/6nz85ri7/+
Q3FchbMzWb3OOyf3vJeJITSjgirwGml19N72GJ9rl/ailUgFTlH6ZO5HKwcK9r5nXG7dCUi1GzyS
LwLRvkDkJTU/9KUdCP/hEjLwpc9yH4vWvF5AiXGZWRpR5KG3rCpQ0vGBM19B4g/dMe/4C+AFsicF
AzVVYs3aJrt4dX3VIsh0i5XN0f9omFTAlAXw3K26+7eH9nUyN/+kPlDya5zmsShRT3LrEwq675XA
+XRke3PLmNh7ElU79wr055gqtPxfz+MHE5MvMmGLHC/p7nOs8GXEqDgliA6whXmDN3az5rKmPrFI
HH4aEK3AIDAglGtxAVUlkF9JkfjfaFAn4FI48uQ+QbSTXSy8uDwrZQc0yn3eaR+M2RhxY5mdcn+d
1hXK6zYWCzesNv/C388KNddVLs8KL6AuOjXlTwizJsoMYlQifpyxg7fv5dF6vQlKfaoqJJGAbgxy
HhxacR02SGZb1SkUwUcrpkmgWpNrwMj07b6/DLefbVPaUcuROtFLZccpYmJGqOdINSpxb9ZC1ttC
ehstwyvySmCJKG0pzShx/L0ruQj4YxMOlFVNxKmdtLivXKFlVnPGruBE6uSCKkNtYyReDhjDCn1M
kRKFsB2NCNYRXTo7MaF26z+mCBIVxajhvoBl7Sit+vHbHUvj73Cvs5EY8V5EZa0Gh7LVHDGiiPPo
l4z4DW6OUrcui2epIO9LkWsHOUIJ8Z2iiq0FXO0zjPxvQR4999jjgZQKPUjUXKcvWu9d+J2Blzi2
Uc/IJMMqIBWXmW1dQg4Rc0gyIRPAw9anZex6GZd9/1d2ocOP/AGjLsukCBKIOsR2L0IKOaMa8NRv
qzJXja1KbCXJAbkuueRUxWp32w35m5ZOeuwK0qbuSUTgm0e9ca0s1A+fpRUhnNmG4URbUeguzWz0
jUvlbLD+PUqbugcZFJ5hIEJ9s5Uq7LKhfeZXrVQ2MmOVMvzA9Y5Dc6CM8Em4JcOzmhhJG3xK1qyB
YhQC3qbnkP9Q5MdiVUZdkP29p4maCCDx6guHZ1JRElxga84wwGeq7LoreF/IEgi5daLwcdgTnyHL
qF5zmCV9ue6UDPOt7Me0pwmIsFoTQhoChVpTwoRi+cV4SZl6Fl5VnSSvI5UaC2+7t0lzOy13ARlW
08mg5/UmzvsV43cNgICmbfj9e8dFAS/1vDGwOTwZmW0li7l3sy70Ju1FklActUoyW8jms0LL2hAJ
PgrOopHThdGD3BjDLyLiCzIeONxR1s1gJxdv9yzMrPVpk6i1vAsv+NCh2U3Zfe2qwcON5PDK0q1r
1SwJZjKViCOzr+pnq3kltlGH8uWtFDsA1UbRJWwPXGhC0XW2wdkCBG+4YM+iviydhTHIZ9Q01T0f
obx8XgOJv2dzHm4ksBsYKIN1EDA4q1q3aDbknUMhs7Sbuna/iBzSv4HI7Cp3OdAjOjKDzIBXvHhN
q2cOofC/5dGov0RGFc6Hqmd2XRlAttY4qIlh/8IVDs4kI2OiXPuF+lrvNx2h3y7kSZeG/ZmYU3bF
v6uxg54p8yn6WOg135nH22en6JBQ39yA91m4ff8CCGpIs4tYw2KikW9DrM1Gfd6aVH8LjWhqdI4V
Lbp6WDP7bBDhI9hgED9+6fdB5FzgCIYgERtvTV8euizQSMkL4TnKuk0MXfSAVJzmmyKyvBLy80s/
qd1EurQvDz9Orn3UuFO6z73mlYIrMqwBsGG7GPvQnfa/yHPLOnh+qYc+WfpLJBrRWhkUBFofPvda
4W1GcvBcR2Q7ix0LFBHvBE3q3BvO7CNqNqabmW6dTrwkeWWIgUcClkfHzBgftaIBN3N0sSLPn/m2
uKZuRV9AxDF5vqpf0O19DdI+7rMH1smP86EkivuT2F9RvEHx5+c7qF7dMdAf5iwXNOrCEs1jFl/a
i70+3XJfx+XkX8WS1coZkkj3W7k5GY/qH0Ukncp5/RfWZnExz/H/WI5zj295hvA+KrnoJBqRAISu
Mr4lMP6apfU8KP337eMHmwWyfz8xUcQiNIVfVzPPCUkka68e6iUzJZV7PmZq1TTCq8kC9rv3fNuS
Pz9iGYYBJyUtYv0c9BOsxiIawIeawooqvp02aL4n0hjdKy+97aJ0q6s8gteG3iJYWRcQOH63eAl1
Vm9J3l53D4M5q4ohct9ZtoTGV9NusxN4IufuLOEFHkjIApW+AFT6aTupWs2acz8CKMTuEp9SJ7WM
fesWbSUDEYCwsi8wz1QgrrM7g6rVgWk+zzIyqIeru3FwM2VCXl/FB7G2RuEoeNt/+kleRGf2Xf8U
UY2SRDBo7hV8lIV4kp3RGx9HbsmoxI3JMf9SnOe14vhWEaSdBqrrJvldTi/Ic/gEbpef5+9+hsbQ
Iu9n7lg+7Vq0LB9w/lFRGfSm4AR/ahuUp3xgyjEPDKLOLIUNRKPX3Dxx+1gGTRJ1R6ufObJEaC60
dbUbIGrtAWwSgJV6A661aBYrojbnsERjUVnuDR0sAIo/nMbRnGrarWONU7Ro0YgicLaHa5uy/o4s
mp38WHOYo5sYguczvfrdcoICTbrmdT2i2z2eUZGBZOCBQrziNQWq3cDi9qhxkhyYoJRRQTSKFj+y
sR3bpMT6cdQRlQQc3bl+RdoJvqegxyNtl7R7zi8GhflbKN/lo3buZYP5vubcmR388gJ2jNvYJnKy
4X4HjtCEduNzB3vtPpRYhGnyWLMljVKqU3lhKMZ66scQRyvt2qKrT3fBpvZsnUorYy/Xsw68g25l
2eqJPzOonlIGtuLU0gEHSWywrdys/04/26K5yizDCygeqxQhlKEfilWcJZlF8zgG9ki2b7a6aVn+
vGaG7Chtvag0gZmjALy06r5aSde/aLBacfcOv97tkxRc/x/fBB6skx3env188UGiSngfarnawDbh
QMZciZLkG3C3GTUU32qQ53VVUYHNoPKTrp8jqwSOlNHkANaoR2jBsQPJPpoZ8d9rocAKGUXtaBOF
BXS7Z4A/F+0BFozMCggmizZiBNMMMtU3x2aWGKpWKDFK5OVII2BUVs0QQuMboqYGK8DvUPD0X26q
ptHmnJLkje6h0P9NR2/weCNioVSmzNzqblrPl4eX/GeLtsgtyiuBYlTYWUuSZxMyU8YvDopKbBUm
e5vmt7Q4FIZ31+dHgXPv3ufMCHNlSY7gLhTrEmdkhsqcATxRr7XKRwQ+FHiXV89PTZXudJais0Xu
ZGAWO++86PKeLBh+kqOFWn2f1Ldz1vA4vGec+3PrMlCkReQQJVDP5qv9EU00wLLX5JCGGIzJg0mJ
rnJ+URHAbdclEnrI1HA9sS9GDCdus7sAG9vJNJq3IuqGgYIFjO4PFXjT7PMisqFMWNDnvY8DuYXa
qoHwGw7FlV3OT53TUHB0dkGljog3EqkD9nyWvEURLFV188LkcLsnzJ1/D7VHWqtEOt3tjFKE54jK
MrSLCKThDPlUs+ilcZM0amCcjgkYnbd3bZ+NpmQ3ctXX+/zCnYZvvk4O6SKny239AP4jSUhLCm4+
NKiBmyvgvZ9m9ywWlIWyAisP8ywO1OG0FGfZFaqzV2zfSTCQWhZ7q7l5nN9zH0Z75UMLVsidmWsW
/ifss1le8abQ/iCdbahmaJ0fOTjf55EnC8U9j/uVCSfROYkz4FdL9fnsCy2PvY6MFnkjIud0CXa8
ZcQ9mi5/IWPGNx6hN28XwiAUCxWrOaov4ZCUYW0gY5jenU+OpU3vNNljkX/SsoAuLc1r83zXhHHe
I6/gATjX7EAiFnujsAZy4DRidsuMbe/Zlli23GRBEJdpN7JfpF1kuyQ00dOMzifXwcBJHVg9G1Zf
Te7tvaafOFoySgAaj4TlrHZh8JN/sUm6aUWO/tXZ1tFk/Ve1s98RkErDDWGJ46iKjcnA3qSWxivD
55RGhuhDcTEYw6nFQMFmZkZip1jwwLjtJc9ZNCguCiVvCJPpymMbVY665m9Vqw8Mh3RDufeYgQol
dqj5ZjGtOMvdUbCa2f3H9jorq6wBy3Jyf4SgRAo0qtYVDtdkwxYAW37VPOOMd7r60DNqUDPHM3CG
U2LBKgKKowOG/aaJSZOXcXrvxdPDvyEXJ/bbFagJEmpXoEm9QUgiVJgGtfFw9D8wao2YQDdYLyKB
mJcHaet1NnrH9HYtEFCgSZyUeRYoDSEzcuwKOoyCgTyjuZvjZEs3JAzH4fHiMzbaBjz1xotC7VtP
zgkvxkrzeMOYBB5oXFvvXp1ET9kYsvxobsUIneVEiIv9qmXTMmUIESUnmlZ+JtAuNB7XZt5E8B/W
xKJqKC5RIlUxS846r4uwz5/CVGeiHx31jYqsO//XyyMdAUq5d980+k5K76rf38bJf7Zs5LwOHvwC
D6NrZvm2XHrKI8Sol5UwISFK9BGxKGDVtk5lL00oMByTtJajUOaB/bCwrd4yVHroAzpnF42VKmjh
cuK47Bi/TYRBYmtuhY6VHiE8qeOG2overcHip3jjliotmxUtvFraDGGNygzLmGKM3BtrPekXitlg
JP2MCheLnpkg+Drqj5eemJx8myFBTQ1xj6cVj6zEacxNTQ37zpL/5xdiMUCaYAPdXRWtCllgePnD
LbLH7BgIKZyANCk878jldSs52b7hort1Kdy5OKF+/bM5L/Ap36smOgz9TBRT6w3k11SUm/ixQvyf
D+7/c+XrDT4QvFgGs/BZiedA62sN7amOgx9WR7eofDyvkw8nYdysQTxPdjUcuHfunXDgNdgTAUIk
ki4Rr6YKRTyjQpJpkPhzHBgxtbWaJU2sJVHwPw27BrYaX8gholnG/6Pu/xkAMh3Hbwrpv9KJzcma
a8LHEMPeTNzBROVcCJ1bCedK4HN0VXIgMYCJcO7+y90h/F4cXRXHv9ImnjN39lrjgNIuiVVZGiHW
7VXMfDp/aw18pyTSgqGQv6Uj7AHD6wfX8rIrD5qFsyDO+1G/ARjQfIkaMtl038uKOzdILfoRaTza
xKpY4cCTSpSfYMfw3HFWZmpT9LRuxmpd6VRnSqCeoReiQUZI1nmRLfRlxXjdclq0BhKDQ7ICq63f
Gb+vnO+tPEnZTB2XzJccbmk7ZG/j75zON0pxyaR3fzXElGAPxveon9vZ8XaiQzMXgrNYPO8GW2F4
p6IUUpxskVKxCnAoDNh/kL9S7cqPGn6mybol72Rw5qlEA5M6nEmePdr3Bhb4XqvDZXlLFp+AQg7j
kz5wZwZWJOwgYllNJvIxPNXYIysH7t3HZU01i0zCRd82OO6uR3BAT9OxyKAM4z16QH2j5BANvA2s
V1k02myFQIybMrOw5/E3nkvNWhAGgOHeDPolZ2Upeww7u0QqerQqQvo2pyHWLB9JaWuxTr0zZ9kd
OWllr9NnoGFTArH+m5pSn3SEfTXh9bH23h4u9eXKv1K4uEtHVmFToyv7Bb8aV8AN+qJYABJQZPmB
gE0Ix8JABOKgDWkAQx3ApTfoS3YkPHwpSGfCrzUUxEn03JEWYtHGdxUY6rR97B3x+WmGtZ0bVmVi
C/FF4OKvWKcIFUBX62f/rHukrUlcDC7VTQ3UW+wIWVy/Zc9eQm5JotFf2QmSbSLOvVO78o/Ve34z
yGtPGivBwuuNMyvYHm/N5Dz2ri3eOr85374kyHpKzwXTqp7yaWlv01RoOSCHPtTV/5hxqYapBchc
5wGtl0u1h7vMD586ck9/SVT7XM3Nxj0G74P+auqs1GH2L911HBUxOT0Sm0WYK1QOQj2bXFPinTm6
63BEisdxCZg09IYtXfD56nApLjjaJ2XyV+XLekSMKSkji1QJN4MuDVvZDdaJTkIgJOC4BqeOPFyv
0aho0/Un4h2mAQYwDc25gNEl3spQRYKhjRNMkHTp6Q3Szejdgze6naBqnwG46Dv/VzKvO4qofHSy
9yRveozSaJu0cUsdGxJG7fUKIFOKgWKT87wl01memYWcvEPu6G9K52u/aPzkf0tUpNd8MHnNWxRz
go2S65LIN5HOOzhlUQnZBcbmuiG+dqUJLpQwNJoBhP+sckWhLshGRQloze2jlTp+iSh68V271wUN
jtmuv8o4ch64txkKMrwd8S39zZu72gCtOsd9Kz6DcjNR2LX5/LKXe9jHKNjdUz0yLZDaSW/tyHJ7
orIsGrSde0WDstbsIYTcDkhjaU9kSv6O8obZ4MLm6mWiTtOBRa5bo+emPY/15VfEElwDnQUC+1rt
8U+rcooQq11t/k2U3UJtcJva8gCaQrrQ6NBXx79xI69IIOj4zDRh0M7s/IOCSsiOBnLBborIWO8p
La4Hg9ZrQSEQY61CNKyDWXLJmyAZdH7SMzirolIwHWd0CLJ9ZfhceOYDnPUdZLYrnbSpRUJ3YR/y
S5PiBYncKZhpwTOPQv6FYeXQVKxN6CBkwkTxC3eBgP+RqbfxSX4VhddWe1gRKUhBFIwFx1Ge+1lP
f6nIiVNPuNS0nJGfZ9K3lmkejqXhWSYs3XK4sg0XekvSFqW9ETkCP6JWox6B6UxR5mpfUhdLU2D5
XRJx3mNsJtbluB1p/3kTpNFl+TsQgcRaYGio4Hz7d5HBnVVPuMRNd+hqPgQtYflhZlxgR3oN5LAY
mOAL63tnfaWbVxVbUeIOmRP8qaIlIZTuoVt1feg1p3wOFBjPjW90Mkrme2CqtBD9atrqt/XwOH/h
+ro0a+hoSg/aFg5ZfFzOnKvsxX4Dl56KAlJAD2TJ1/nyJ9/kKZxAPgR4hyWScO+6eBYYD+fE6910
BHWXwHdtO2et1QCzjV1AC/s5V7gnS4CFnvk/tbfqAGZQfBDCwR5hGBdDhobcfuh1Q377+pQMzdtq
96DYSNl+TFvB2JIqeHnOAN6kHSI8bHxkqM5RS4/qDZ5gKePg4YCNi4Vc0T/ET7nXLoz566vDC1az
cz5vJ0SdTYlQaWOzia9cOJGcYgr5BUXHi5XSc7IAPlVU5nCiCqk0fw5IuEObTATju9FT7GZQXZDE
hPm3e4P8pbUew7KwneWQEN2b00J44bUCUGnYDP1v+iDzZA80rJ2M1NHYgUSE+i1gSLS3i5nsuMCc
Tf3z5nSwpcS33z70JAutkd14vYfv6rC7Q4dFFbKlTpFaPKXHWthFtyI4wLDxMnWVQjv2d035bTzH
Mte3PahD5tZRW2rM4daAGGYbTY/Gc+paL43s6OQ/7+jmB2beEAmOZWPadH9XqaW7lOt/eZ0n/POo
uKvRi9MiA3jP27EerEpazdngrUOX8wYoij9TkmJjv9iNleibnl+esuH5I8RcU/XbAYmnukjVeuGB
/BGaKD9tdKgwuh8vzYefTzOHEok1B8vsSX3eOXd26HMn2qw2XJ5ZfEIw2Qbr5+I4QMGIbZpDLmV0
/a5+syHK+sbEX8Pz5jY6rAxFdZ0pR/C2CAXL5b3Fq3Ve14zb8pJus/CyWPRkmnPLKY4xQQhjJVNC
eYul2EIzog/058LbVOWpF6wJdw7NlwuPo7alQ9aBWTXqMh233lfTDMGoEnqSaOA5v/K5uBPug6OE
dPYKdEw7aIiJ5cvFaxzwJKlVyqa7VQyY5J14ciKvvJgZVojM5HiSDtPBo6Wo62Q8x7t0S8lUQY1w
rMV6Jyvh+N2qECdv2uEvjOajun9CnUFsJcGfH42WfHIAmwt6D75cqhtU3WEZv8UxZf7w/gnMyAqS
DBt9sKJjzLbFMEGRXsYDviQ5VjLo+2Qfx98oYc66nHwlw8gHgMwlOY4l7fyciriezK06BL7mQETS
seCZztA2V1SqBsn6c3qiKMsoy3EjP0GVheHF+Z+fVq7F5tvWoUZD/0kt5RE4j6Xzdxr6XgsxrrBc
ki7dJQo+A+Nf595wuR0VOaofREQbrY6ea4gxEeQ2U7vCJtdL0hporEm4UR6a2W2HTb+q6ay2cV3/
N9DeQjMaU+RYCSAOnNGeQzcC7icYxi+joMsPzrhUSRdJXsVADiMazAEF6sqc54On9xoSHZM0ahKH
hViReIZx8hScb5IGIn1VEYw9Aa6ia5NGvVhJXxKvRLe2cyVGwlUrDgt3OkXXw4L4c53ahx9Ivjup
ev22ea9D8MJQ/F+Qg8CMscyKHeFm00HGg7v5qniIWEMvDLN0nsgCkjK+NCzu8Rnq27/o23161/xD
OPqHNoOPJU3L77ORniD7fEGsj9cqDvelfSfyta+4Az/raXtmy0/RfaPuUCTEaRZZyRRMA3VNIsuE
GwlpFZIvhuluTvYfwwzD2IB+XuFlxBy02xMAEJ5PDvcS905dzoAIUkfLPw/CoppZ/x9tvxDpIYMd
rUiYPb9I5Kex0xaWqk6DLNWbxHU7Lc8muU+JlE6bQDXvdcuCA0ineWT2rMt8dxem88vEwx5V7nhj
vzYumxr8+B/tQpx982bVd3UbmxKaVUaz7x6kc8sUpmQCspzzOxOUU0BV2MZRK+zUsdrwC+OMtP6H
jGOkmBW8gp03WMkanvMEKijSHn6dLgjiQ4qdqXStX6ubiaGSP268yAn8rNrwkNlPb7Ux7AICnUN/
AXCDWRufnx9FqbeG8B4D87GYlCyL+WT+bsifXHdspcA/s15KEEsSgnTxp1gc8141BTbG6aeUVi6k
oifBGwkkoJf5VGD/0pS/j94/Q6LSTT3aA7d0WtF7RQLRJi7yWQS0yPI1/C68+6iJFz9ULHyL//AN
Kpz5FXP2gLTfs4ENQhMH+uCOk6VkCVziv22fgpigDEhFRT8ik7ds5rYjSFz0LnxKJnY8m1Om+kmX
+mFBC9wq4dWUXUJEEYJ19S8mn3Fno4l6Y8CHkftzl/YKsOsZ8L20dbLFm3ZQPjzXuVNB4ATWY6bC
qZAN68eRSfafhNxqqI3+xnrgyDckgkqx36wPtye608HuDOAXYPFYTNCOwO2TNCJXbbkBKZigK7jS
e8lXm6tHO3SJ1oM4ypPqAp7IYs08d6UUy4Af5qR35U8dfGEJ/J0G5wVCMx0fTz9D029FrqLDa13G
E+nwe+/Tq65cqGx30KkjSJ5lXrIniSTOgiZtZ2GQwpuqfxWp/j18zjJklvIhxpJlwS+3SqH/PIe9
GAx/hNvWCd+iurKiDlgPFelV0o5wDhLLIA5Fxd5CivXth6fmNpAyo1GFMv+YipQiMfRKB454tOs6
x0zPHHkOEIxoCgwdkrcMpAhC+2SMn1lOkoBYDtJt5E2oGCE8L09aTyk4Zg0zZV7ys8t7JQ2VEw/8
ce20NPo5mtPwnvWTn3MDkfrt7lPgfpUxS6pzHllZ5yq7apY+ADKaMJQkpfcSwb9cq49012TOxHwT
AJMVY/i9JFpWNKEwPgAkx0H7NTi5hJYaI6tHBppFI9a8XY/JYOWiU5koZ59u3eyTKgJbUdqUg4S1
Rt/GUf/VW0QhoXj0z0QZmDiM+RogW5gpIoQlCU6vhsFIohT0YistUWx1v39OKqk8lMdYVrEntTHt
1RQ+vS6AHr6v+2CL+hd6neI6s0z+hvAJcoJrMCYK4VbgPdR/YlGhy3p7/zY58UQlm1IaXFWXN41H
Io9uuiSInX6dkA1BDvSD+8JCqdqEctj/P/OKG/DFBspfU2NFVp8jZBY3ocfxQRgnIl8ztt7+ipKH
A3NiCciU6pUlPhSU7YvxQViyXNb806AhS4q/l0Ik+LX2iNzmqcECtrPkhtqYdY/9yvCvARwxgLA9
5f4IvBTyxkDVUX5yfo01pBNT4Je1fy6S8O2sAYsyMJRJgeA0w85UbaPrqOjqHhqNbTenWb+rUIBB
20H8eYTB57dYgmO3xICd+kNNZglGPvJ/SCy/bcnvrbTZfOmg15G7m0jKspCi/zgEFFAadpy5YJ7Z
YN12XFn6+gK3+xnzMlYxoCxoYOJaSlBHNX0hqF3HDMr4Mh2IjUqEX+KnNu6S6GoaZv9LoFGqJR8U
kIt4bIXoUsbX35vXq+WIurRk6f2DdxW2og8wETKhJ0Hvh2jbKByd/M4Onap3FdSsd9mia9k+Yil4
vL4kdgV/7C3Tf+BjcOGHnGqB/5FiOkK8DM/YpxPc7DDjIm1B9+kx77tLL2hrR68hy3aKWjy7fC+U
PPb1rO7iLM+DyHlUwYTuYMQ5kFMzSxrGDOdQgv56RL69qnpuiJSX7ntr0dHlEAL5p3+Xw5kwNnpz
9F4wcLAJODWbDMSPbn184jjaW2RuBPI2lLsdLPU63R/557ib8NymPuUyqOYHeftj8G+JAEIHlviv
+vLgIfZIRBhgy8RFdg1ctuCLoVURzh2X0X6bHfa5cF0Gzngin9TKmdOtoYa0ahFexhv4NgwWwt0v
CnZQJ3MbY60lKkTM18+yDDvDdYE4RWeBf08WoirsovLPSTzP+GkfkXabBb9fIXy6p5RoxGlEVd9b
hM1w5iGYc3ZUEhK7eRoIK3cDzhNwqRGdeJyo23X5tRUku/QCnmalVskfq8lnMm52WgEWwJ/N3N43
tggQX3ctrio8hlzxMGSqf1U8ykEJk93vlcXIaUs8x8TsmZBJqyGOeVMh/NRjxGw+AGVxXFdvjbWk
5FEi5CE6+jUyVMVUrk6smGTONLW8qHmLFS++fovv1eRUQq9rZy12oqKB4RFmNf7ndCPZIz/7g2eN
brtxfui9B/SuI0IBnjYrRB1RZuS8foyhbs5F/hvLE2suZNwc71+FSATZKy6+93AmZ2cmzGgkz/Rd
HoroX0KkDsFI7uC0NGzMqqDns/zeNLeq67qjOspICfWFximMczUYEiEPFSJJl+GL7HwaTRgVt42Z
nwt2WuLBgIomFsE4AnMrVtYvcJuqeRTTWC1DZkzmowX+qMZAFCUu5QWx/gfS/jjJ9CJ8iDMygOqX
bdkKCbz3QH3W2zSVn0Y00btqM7ufUSPyAVZtDU1f5ELVRYxbwKYU90bRN0iyOufaEvjLNppbQ/Yn
M1B8tiAVxE2oQg2+EVRLkw1N/Yynr8p0PhblRN0r2MyPU+RXp2XuM5sNJeQluZEAuJV+ZoEP2cZV
A9AnvPmPHvFv+dv6ZgRdqM6l1PdPB5jIB/g6h2ymCaVK4WWTgQL0FPuiIm5IQ3hfnjJwqzljzGpo
XqvIbLd2/hER8mV+nAtPUITwTbkKS36G19ImBM9spKAb0l9jaO7bk8SR+Ln21p5H8YgMj+sgovOp
6LNADwhwmyNH+7mUbPj0hiXErqYeyVfA+j7eWvWfAyIK5zbLDjqOG0NwYjPPjJF+SNEGYZhrM+yi
6a2QSjrtuKEoIxyx9NCY0i6z11slztiRN70JQxYwZuBRKYuVBu8FaTqlC7APzO6sRlodRYevgqcx
9M3QH5phvAaWkhAHAywSV5C/uw0lpSgKQsOWOU9NT/gsNvDdJ1X5p14veVDQ1uy6VWOc2UolUoz5
jZbjjFGHMGJhKSwJpTP1J0t6s+UXfoy9qWRENHTMMrOloybl+0qYtMLCHNuocnwK+b9kQA05GpW5
kRg8qaaNGZyF+Q7aY06YoEHOa6xFG23NGPGEedcAlwrzlxkEn3BOfgS0b4QypE9aM55l2SZKw/3f
vxlA/e/3bJ6ForcRabKjOmEWyTAJNTQmjtCEYTLdvKWhh/5moudTjeijUEAMPOLjakrDyH5/Ho31
DtV+CRAoNR4XPjyfHcgr9Fc+XT/RpTn83t6PgE3gse7XSX1oY/WB99CnY/PmDFz8oqoEp1Cg5aAk
TWMpYrrG/NnjEYrIVLf/HXzXpVxdRwQ76Flj52aGtZ+3ydBrNLRdb+dbAW7lZao+WPQ5HLkp1IY+
ajkAgkEK0x7neBm2IKrsXO59uKJgAuhOe8dZoHpylD6I/MW9BNXM89XAlNWpv7+W6OuZOlL63OWO
dMZcfqP93HTKNjJMD2/rWQemWX6WX2uqxHgFQe2lML8Oc/vxYkgQSxQaTgjIdJF0k9Qezo/tbuim
CT0ye/QVcHR6xVj798kOevNaTaVDET4H3u6kX10tfFiZKNgpCzLK61qAWNkRu3ffgrC7kLIHhI8u
GLPRxCV7nu8HOXbwZDt21Th2JUH76z3KoKDvHNjQ/SYTofM9uvYPIj7ZaLKCp0EXbC3NIQBsrE6I
aAmVH/Qn5pe5zT2VQrZDzsPDTqtcKmPW0jYZjU+IxessJfGuTZHi8oSKZQp5VJ8sm3e7g+XdpuVP
7N/pAW+Y+ftHvjxwfP1hfH/QuvuiMqsrL5SOYmR0MyyZEa4WgoS1y2Dxh1p0NuL1TmFJoSQl6hMP
QBwSe6F7Hem3xuWljhV4ze+ucsp77XKOZmDgGTSd/9GW/bjhC0sLR/EDFNYUnAdiiG0MUNjFmDmp
Ii0yeamILr0I4zlj7oWsUDCjkUyIOCvTyUqSTAK0MhYGePpQpSgcTVYyXpZpC+9P+kH1dqJLF+Gv
sd4GwlqVMzyMar0ahfjuNXb5Tz5+Re3DnMbYF3B+JU6ydSnzX0Xsvodk2v1jbS81P7TEglYlVu1h
KbtfqMqUbPwdI/hBDrHtCztepT/iPy4gyqZXG9yUqIQQTSaEkfocrAXI4HcFWG4MgQYUmCe/3cTo
S9dqmnCHNdjRQ3mc8ItOULNJ6a+5oSkQoaAifBD+OZtmbne8AkGCi0yxGFAlH/mdzKAdI3MdcM7x
HTOcjPxCwacX/o+WOOjsHIg08wjUj8GX35DXkyK8q+b4uoOc4N3dwVI64IuIrQlCBgktBk/qv/+b
N+yRuzkaMFEjMXfzdNH8k85MDD0Ze7KT5CnerIzJbL18Azj3yUEq6/WhFnJf7JnCJkeMvhPFK/Lw
iAFA08/9r9X+JxJVXXJy7d/3bmZZ8dspimoozpIYlVSdmu6LD6N1gr4Y7VqTvRoJb4qnclrGGgkH
3PMjMNWfCmdjxH2JmP9B9DlF6up7A6ExdvqdsPKwo0i1XGeRPCUcmKF5/qPxKx7kdxcEaNzrVwoG
hYXnigfug1rfxS5SIBPxtHN9DzoRrE8N1Oq2jYuicOSZ6ZQwP9tMRGjZio4L0MnnVpU6wl6GmrZH
hwmNbur8ETaCSgpaRgSKjVnLKdVacML/cl08oYrFwl1WyirJ+Cog3VXEzMb/JhGQEkUyGTp73hKV
GQU2QAPJOyUn2sYVgpv2KmOEa0Wu6nxpXFt0w2H0D7AKTLwb6u9Jg4ZGvl0xgHWB2Kil2HG8xiLe
2ORGcJc3Pkkj+yCRnO1ekqi/M7GVjwh+5FVNHGfmNs6e9cSZEmWG7e8SYjDU8SlTJCQdyaNV6j24
1axOKngKsWtpUPvDJoDj6j4wPthshDehzweirtBzh+uurOesXBU16oCwhG+2rS5rxqcwX84yXsUU
iTVgp5KwzZwAz4a2bKzZEaznXbv3Dv1mH+kIFeGi4JmCkJiyO+drp1FvYh+G2rmzvOs/pe9yiodD
L5dFpw/cKXYSope7z52FBhXC/2hvIzS5n+IGr1d6mVGm3I2oRKq8lfHJlhoIUAxXlhpkB3myFa4l
odgNEg2cW3uJ02OrBPd0UG5LW2lszWDQvAuH0RUnSrRBLolPGlLXqfIli6od0Sqnc7r7A4J+Ipxo
1J1r8lVicDr5LpULrQhqA3qeU5Oa1Zzj0zq20j6IRtHkZKuKTx6MERx+idszARm5HRD2AIRkZaJT
sdUU1Nn5JxU22JA6uqbFscfgZiLZTAMwvL6qIjHduQQCThd4SWxgLv9zNlFH7AykcygkhIpTEBmN
mWn68UWK7ACWsxCEOQq+WBOTD25/41VpL+Vj1sZ92YG9hTBEb05HcpJd6FBRMIb+95U9XGad9Kkn
5pUL5cvkb3lgMkQ2yYflFDVdDP0kb7p7iVozN0k+gaOkilbPynsv4fSViezU4LOH6xFPNw/X3IBZ
6BvtUsUnzvRpTD/9ab02LJByfy52E2LGHapupTjzmshFcZTTUohZFxyf2qCJA3TTtcf6VJCWQdP8
MHZ0XdXBQBRfXXTVP37uD+5w63Kya/rkfnb4U4Z+677kl7XyZ1JGxeceY4l4infwrmtONJ6UB+3O
luGEo/pbiV6GpdHs04q4tXmmheL/M5iayJLi9rTyaElD3dWSpxBKC6rQ69YjQCh5dK/+Hv2+/Ln+
S6mSI5i3p3gcbH29WJ6HhpPUflq0r2xxGALqwvanccRoH2p6ip0Bef8ULbWhlUncW71Yn5nzp2En
+R5gki6e08cs8ZqQEZyTa7soxdFmYosbL7MazFaX9gVchguh20H3BhG8j48OIea8E1yELF3POVMh
VkU6glFipzQ+dBDLp7wTF4NFC5S8W4Cr5vpLTLq+M0Ro7wfq3g/vjXshljiOVyG5GBZfIv2gJ+V7
BKgdQRP3seOTQXpzebmR45ZfVOb1QXTnKc11FPzfOWa+BHdL9AiFGttRn3SCrX2GXH5hm0fFPeLS
mCRLfW/tcNP/vNCsFOR1V1PzMrMbv/WU+4MpGkyHctLqf81iNKRIUaOUxaAnYj6ssUy8u5vHcufu
1WMzN1V8p/OpSJjpWWbAtdIkLIpNBjmtMdrI/tqZzaNu88Ri4aKuawq7XfzC7x89S9h3LdVTDa65
A1wTIHoxfANdS10Lv9MK9iz995twg+EgxpKSRMnwAeCINSU8GrX2KhPWSg13fOzXm6Czcfw7Rtx2
pR3gSfvAe/bChKHL4+weubNdDrv+w82jtZz6v26kQ9vJFjOGjj1/h9cbRnXyh+hqHFUA0u370Fma
L5l1JGtFlRi5QJ3G3la0sZw+gSJFT9tQYOyLI90LwFDqfhs8ZlErkC92Es5pDDl/Y2Adz3pyz+MT
heoPcbgSDguPAW//roCPe8/g34M0iBHDVOJsbApi/+frQYpAvM72ChsLIVd7RdDnoPn2lSd4yu1q
PiUPpbINwPxfLJrFyLdq/48kRMW0VT/Upi6n07osPj23b55sdH4mR9chZQN5ACem8QgEYORJa73G
8XVAVPSm0XoxC9WusIuNdDvAId9E6IwNhV02joi7zcPtfzXPcDzhNdp6aC7c/nBrW7f8/OMn8fTr
8YHavRQGlI1ZNCa6hTTKa75b8gZZdOOM0N9UoKtyRTAhNyYVvKKGMwdT7YOQTEvGQ5ByTCRCq+rR
lZ6XggrmyxJ6PTFDkQ9UFCh/RGrCcp/8wouGecIx1wLeOYO+7eT/GfZYtUDaSRS/rWneuDrF3fWY
8rU4PJNVLzMVmaN4LbOIkGZ28U4ZK3TuBR93Qsg9XGvi6z5PQw21VWYcd6+EXvmeHxPFwqP+BQ7L
lAym9A6aPAmsG7qMjT/hvT16uvezN5YTkFP6j/yH9mhWBBCl1dfUr5fVoxj8ZpyXck1pCNsWOul2
eQewUo6wgEPIaHkjwrpd67WFEaUnIhAYvspQKMhYdjRm5SAHTR2zaSpa1qAUM4zvFyQ1SzLyWHIe
lm38AzB8s64VQnD1zUcwG7Q2xMw7r0fzKHuUUF32x/BNF6mGkyuBTzvDzZcaXsWf1Wn8eLjmUcLr
9s1TWDaNiIsZBycxidr8aHJIre4Z03uq2TfrXym9OKDKpB1u6st7H0N25rV2aIQt6P9zkVM6eHpM
U+I9CGODMVGo2EMac7C2h1XVRO63289OCVOqCWINYeBFysTuntLRvc+PpHU4aqKlpGQc7VMweUor
XycR+R8+C39mZs8+eVP6CG+uT3dl6x54AJRSzuN4Z0asVxR7QMCGYvOGhCV4KgVCRchcwwVukegp
aFPupC4002ebCiUGxRKE2uaN6BDIxOubX/vCn75ifhajjd0AlEtcSEB08Ddjo0yqvbLgPnFuj28V
sSUmB3nARjvV6PiqJ2vfXNXs2HbZufO0A+eXT9BdBP4dYrwlFnhC8++OJX6r0FWinaqtTiLXp8M1
EQn/oW8SuR9sBxz/ABEju+WPRupzYkcmyPl48fFep1Tss0dhWJ32bsX6KSaVPYN0K5oWRpyUhx3q
TB3N0K73B9z/OyDxN0wglM24C10Epr9OqtCxjKz21yt9oLa1qh+iIJjY0Y+rRDOiFcVNvfhnrOld
Ly/yRoKOTtJ7Ciwyg3pSK1DvHruPW+pjypNRV0MX1BYmFb8icoOqqYGTlJUoSToUIQdOFUOMDsGw
PxMuVZpV6nGb61hBVDJHuHJjNf5vKzPTzG5j2u7pUbUwjjfeYX8wGhew9Z4D1IZP07OiCW/McOfS
v/e3J74VfdmGjrWckMstn9etxbIggNktxMYFbsVD1Odspi+b/ciEosMS47LioVCUhNqgFonRoOAv
Re35GytFdZ+Lsu+ptWtr+zjt+Au5NuL9fAnbBobDwc6ElvN2/IivzrtNNiRLHpAQygxYJUx7quyi
C+eFiQpulMrSUvUVyQrPBI+1bwGwDnnyWdvSj2d1PE2ktDhDpFHMV/U5nA2S2sAJOHJuuuDXlrdO
zIX+PeZHBawkmtQptjkhuHOvFu6LtwFV7Qp+ugcRIQbHi894czxc2YLiHspXNXAGY09/7kG5zlUM
Yn9JlDb7FbjO8bhOqxyrII94sfqFUXhlVCm/mcWjQ55wbbxe9SFBiLenB6K9E11fbMgD0j5pi+/h
JU/b5aZtxpybOy6XGUsqYh5BjhwD+mXB//xE+sdlQmeiAGVwoFPdwoN9UlJhYYnnNMVJ+Zsp+ee3
bDCLIqNt5MPeN6CobpsOEzDME+jJSOPaA4O6LHpKqkTS8bpm0RdPqMj5Gz53AmLZfQbnHSgPCNSB
aQgbZfNxgB8v68IqZhjq+hpKZJDuYW9pprM/p6POcaAwSltupO2H3fF9q8BxlUBdIB55FR9m/vwA
iU5/VRcRlsqP4ztyziMQMAQJPPoXd4GDp79bIW8ghWUPA4sIDM5tIm3dTDtw+PVRfzv3VoAe9uFi
ETHmDFUz6XAUI+hRwOshjW//NrGg/4Q3qo2O5mqTTkaOGy4iWPRXnJXTdwnQw9FMjzxwhhUZI8pY
wHGuh3de7VDdFWqymJ3MPr4wOMYGH9SrsJ8yW+QqDM7ECVwjiERS6c4G6dYm3qQPTqn5Uoza0bH+
AB7zdLCyia3ruOUwr9yTWI7aaaYOQWYl8GXCDO97L/pgWMVgDHYYnvIr1Gi+gsgHCHQJITOSJCLr
eCQvNLt3wFLpoeVxxjYEa0o16ZXhRfmHiuJXW01oU/LN19/M3VzY6AdusVs3BxQYcixh9cw+ydYD
k4jFw2ZjqTgncLB555pXlUja2nr9DewW2j02vIlGZ0FbD9KIQtYt87H2j20GYsn/9o8IANhIri/1
ULAfHbJ3O4YUpr+bnAenxFgJBTvOX5X46aaDof3ZK7EEc/wK/z1zY1PjuAZD0roNqTHeuE9f8Ini
h+rZoTZ8wMRqubGo98yfJzCWTzP89j2CrLbpxUqdmwEHHiJypUDsMuHiTQHjAAmN0L3c+MeLXeNh
iuNbAohWeYBT34KNdKUbrsMCUiOPPpwCxoBW8C2bS4x6oQaKP9QCCIqtUAptkFr1A7tGjWWmPg2G
3KGJRVLWSbFyw/g9cohh2g2el3stncSYdZn+9VCz150OmnhmERizR1d2w6zUrFeW3JuHWpfcwMfg
gWGQo1X/DOmsq8LSeYYe/CuuWonPmFNtK4lnYnuPHsRP9A61108fw1sRdF+otXBhaOvYLjhCrTqu
jGpj0LjEaHD9OIQ2VEu12iQl6tHhc6qLgK9Xx2JQeOP0pDaM/m8imwyxWqvy+d78HLcI2tw91EXH
v9GT853xu5kwVq8rB6p9iW6SzvyQgflIDqy+s43nom30R+jaupuv1b5CVTmRLmQFuyM9XpAgGBH6
weuLy8yOmoYcFA0immZUPutEl4zMUSwjtL7i4wlcVhaBtgaz9IKm8q8NSHtPU7ltGeaMQtonRLMq
GnaXY/E/XOqf/WsqF8h/tHN6VwVF1eCvsUK/zSfBbcjMD44uj9THflZX79+yEv7+nFs2XjD2nAch
ajsMBT7bqf4D4u/02ECWt5SaB2sCheeHcQ8T4YIsMprxF5hsGNCf1Q02LBoin50I3szSdSsplYFy
y8biFjNgzEVURu5KRd7xNJLIESIVOFRjG9iESr+D/IadaPLKiNBGEeS/C+CTR02AUpNKdcV5VTBE
Nm5yL6d6Pu4l3/ziay+Wbpg8HNXKB+4A5SLka2cTjGRzOcbT66p1vDsiXGAf+G4R6eqqcQxYd8g9
mJ9KIEMqTSSTC7lEglvw5+2V0QbAY3HIV/lMCkAzWs2R4ULahWfuIPkanlw7mnEKScIMuPsIuNyn
SLg+ZBfTVGT/lLeaqq8iemhQoGr7g5kGy6JGN80LYOvsA+XNrqRJAimjKj1DRbRQ86axX7UvhKRf
BCkEj5j/cdmsr2yGuoIjK2bRa6uAzTqd3Jdw+e8G+NGOsRr2Uzmg5J5gdAZPluwYDtmS+3HSW76f
K6WH9brjH+hfICX5BaotCloW1T0FcXwZEvYkZ5h8mQz6xKju7kEXfJ6QVB2fUGG8+vZYdqo9mIhu
J+nIO0WirwDPreUyybxX2fPzvLP7FWPIYpgOuVcUCsN0sE4l7ZMrCj0qx8cjdMnKd6+vJ1xjpHS/
6bNk4LIWYZZ/6ox67xUcUTFrX2YZseYBc+tMtsF7QzRqHSRqpfbrwoLAX1JTssf3at63bxP7kYH4
ux+fzqDpRMdL2QZjOeB1H6fL0K1lTJBjQ1MNDbCyu97bErYWqiDgCD3N013IZm3Zh3EexDKL0NSx
zuHkl+86T7MoJGU57H0bh5KXL6di0EikSebbFTOaW/gbQHtREfT5ls9qZ3egQLUwNXOHwdFpcYDl
CqBnWozyuL1+SKNjusVCWIa1lf3/T3suq+B0h5AtzDkQRc3MWcSaQCFkVgDyndnHm4qJ+NcbbDe4
FEMXQXhlOaffuffDP3E2Wi1RBDY2xR3MbKD1+tAl5S7w9ZeM2OGoe6BRdb2bZv1fhiebLXPWkigG
rV+KUY7fJPEwKT8TqaPubR5cBx49omfv9WLmO+kJjae/wixyrgxP0H9bPfwVE+VoFNQ0WZU6c8Ne
kBSkEdicGPanAOHiw18/k4aMb4aGDBRW15agETNEtXX68D7n2ZgNvLY32oTuOMutUILMoTg2JQYL
1j1YQsDe85PpntKA7P4rAD4ruuh/znDcDHP11FbmzIEKBLV1gUMp7FT8w7fyj4XlqL8MpKrdzHUr
QlP+hbt+pgzxGrxoHxpDoFoCcXACC/R4/8/4JsMSzQ1FGLCHgQz2GMaobOQnXdh+r6kwG346Mcmn
K/QrpEgaTkphzjtuy7+gxuVDiBB8/GvClTYX9gLvqiKBphvZShInv2hjRdl73jRZtgDVwaD9lyum
obExJXxwR7oRhNfNvFJ0AM/66q20Tmti4rAOOX1v/jTSqd3RQsyAwaApBkMlSVc/o9rSjkVpw80x
NpXbUUXPWNYnMg7bwe+wi2wQ5TTpRvuAoVXU7JV0PLONBLsDUhJfY+iDsDmkxD2tN1S7XfvWobrg
9oJqrgzXXAcXGKXjI2QPxocfY/8h+XknHqaoPa3MdBgxOYziHZUkcnKmlx7G46umS/ttIwLeD1K/
3tsvVtgjnltxJyYzUFqHUGTmjzyT7bDBLBVnQ+bSuADN/bO6rjhi5azM+pG6DLxSyxwQsPj+rZJy
1Rcxy1Uw7IMMCeLKtYpnzoyVerPq21bN9ryMqY3gHjAqnRVd4J8DyGd1XjNA4yuSXvSW+pIiVRLE
oNh8KOn0DJsTR5Vo/FcQ7Q//d7PONenKm8si7autRJ3NweJNQEbAJS0ckhz4RLx0cAt9WHRdXQ4N
Nxl1ZT6pyYrGx1cpcyubXjkebdjlWBjS95u/JBFfqt0H5Wk0Jr+McRFeW+tFK+wvC6B1kLhH75DL
zU5h2NFuUFnZQWQZpKiB2GOmGrvz0c8BX8ter8SVcw3wbtr2MxjTa+LfjoyWvpyk81F0ulYEmNI4
r6CSJVdNGQrYU2GJRCHnm4Y2Spnqu+1qP0Zl8+xJ/VCM4EltIBzr4pJdeU9rCUur+Ff7ua7sSt2p
fP/9N+cHFCIg9e8UBZfW/VNSREbecRlE1LDAZbY8nFHTY+wBiPNYH8JbU8/ztxnD2WZgJb5x90tU
Hz+ljos1H/41WCKNJ2olfUwCBf1ubilwBi+z2B8Zkzy7w8Zci9kgEf3ojcWPALYXgX0yMkxA4S0C
hTk9PC5PNN5pLQ1yt8OShUuFGvsPm7PSEv9uoVDvKpbwdXsNRPgCeVN17Y1M7woeKfFRsn58tyiV
RJgBD0JF0MiRCIKIaoUa6JMZUpOeQV4HvNyJud60MeuzOCtC2na3hzl/TCn9VLNl3H1I57pVVdwF
Ut3HWDJhUOM6PEkn1sX3ioVgNIRuG4VMp97GPCajvBt0OWvy1vCKsxfBziOuJo1O6bPgCBi55Xsw
N/XrvRzYCFaixG3u+MWvAW1HQsyJtLU/BL45NU7j2YSKeYbOxsf/NaY5Nd6Se/nFkbOTTQT37aAc
XWddVt1kt5oWzik+6aCxq079u3jl1xYIAwUFsgoWEOUiPy7txVf1jC4v4hSjPOaNY4QDPdeDO7Tr
ueRG3ScoAH4QXuMnFaRTuFRE0TnTxzQ8lsV54GmdSYl4GNZ02L+i++knOrVuXCrHdADyQnh7nzxO
r4gOSJSxWf31pdQGyfQNsuSvAS2K90A4vF8DFyspPdY1l7JOFF26JLmdbSAvHhnsZXHErFXWYfgz
rgodPWd5wsaOUQbgSjAhz/6M/EEkUDjja2r+JRhCcPOjT95K4ZEk2dCLuO93FyZMF5Q9ZIBbj+Zs
uFOXegUjrxSv/zVzYlTdniJEmypVA2OEFLxAHd3HBMoSUCEt3QsCWutV8OL0YkPPnixwoAV7aPWB
xzZ8eNCRrQdB0Yeq9ZfNPC7LWJzZD0qCL2wU1otylOD0M7xSbOQDQxu+15UEToYTOfr0S+eHrLge
JuQ0XG/gFCJYzOr0jjPPB1OX1g0yUBrSzllxXbrrEpe1tx7+XIR3hWBPExYVd7Vs9sMcFRgRpwOl
re+RIgawL87V2YPCZ3dus6pi7uESxyP/J/bRhb22LvdJtgEnUWFtAIYaGicSX6j5F9l2EeIr3dcF
+8br9t4tQ+r7aQ4XXfxT7bWIMRAJ1YFtkCtoLMyBoNVXvm+hxrPIRBC+cZ7sawDVY7BXoJihToGp
zXwyXdDkIWIVUhXc83HC4vNtGbusiZxoAJV5hxoPOQOvxYfXbkiBqNAoOeGb6yHIFS+9CN+q6JF2
+DROg++EzRzr+KNpnqHsUGBNdifcfNMJSrhjXRKRmptv8dYs3CjYbdgNOluEEhR5moLhl1yFpGcy
oeJ0ldNFEjUPf36YgsQVyCTmWvNXXTUQYfKRgNV31ygrV8qxw9acHpMAsglKbK+EI28G6jq94AN2
r5mV/FPgBirb4G8TkjUR2m1hrBfWlJpUycwIBhTiHFHCS41GXMYnvWt0VSfwNGc5MGELvFG/J8dI
ODRgJ93qBupBImwraX0FLMHpmg6U22NMdRPsXdTtzQL032wSvUByWuOiYNICZHVc6iQK4+1kfieI
ylIeqwClWkY2Dwog+v7kY983hQUNbvLiw3HtYzNPc/By/VyxRHn1XBTk3KC7A7YPo6GKqe/UH126
mZEDfwazjbRpQqKNMGaSHsBhbRWDX2M4pLjCTWJaJv3pT4QSTMcLMuG5YeIUgGp9FvQ7ejWMEcLn
44kMru7s7pwtgRZusG8e3mAIaLJrZGrkhnzRd+Jgw2KtZw94RF+T59HtVa5VJOoZVuoc196V39/m
a2vD8QJuXdEx3pG+cgP9yfQqldM4YctcsmYpfS9ecrX/TICaOTZbBle+yAlXtCRCv54dsej2e6VJ
mdUoyJS4uNTOZTQxG2gDszbQXonOsWXE7hM26msq4pJd6RpgpDhQfpe6sVigYE1pB8l6es/SkMJG
tc4/41Z25V2VwBpVeuZZzdtg7KwTlXpg7i/nIAxkzOeaCyUbzYSitQycqu+lndAyiT9autZ1MIs3
raTDG+dketgYDMVrdfl2W7tRzl0WCxG7mrKRk1LRu36x2Ciw7ECICu6q+BUXP5VlTy7irQBI+bI/
hupMylQA5AAxWRSQdE15FSfTPbQY0B+yzMAVnPhvJvgvTr4Y+qoQiftNxeTFzoQ6tuEL0K1mbw8V
4v23QFfegIzXrHlwXnIjNKoDBDBqY65m/Z95DK5Zt49xEeAnUg82pU6WRtmQKd/DqIg8iwEDBHkn
u9IJwYqQUUhcDXumoo9jW/SdjTSuaSnL7bPqzYfcKuTH8IUwoKIZ/DmEBDJx0k/1gqp1939VRNMc
cAPrdrr2L+/SggobFwndMGormAJqQcPH2zomn2ZwfRCkRM4XTSHbkh0b8nzLg7era/ZFwhNvV1q1
twxpEmfDWrBpEDQPEUHwHUi0lpKv3/7aAaeEIbjCuhZD5ifOXcmJ+vcRvSsJZsrVWjiUTVMTmNdV
e61UppQ+io57LhmRd0PvS2YVVEcigKKbJdqobYPudYHlULLUZ7w2JgYDcoZOV82xG3rjSA9e8JHe
t4YAECs2fLU8lDYnPyY8Ssjv/QxEubSauh1m0cv71Y3Vi7ntq0Y+8U78T4ppVk9k8YkdfalGfYJC
RdLWgutj7bFW8l4u7P7Q38y+gzfuGwtU9m+Adc71HCh7xR+KOqCi60d4+LR3ZefqVng72JjFmg5R
1k2UVZfiJ1XTnCeNPUtiJhEO4lHhX3RbEzh/YIjEhy+n0wNdY48lymVn9Imf8Ut6PHwDDVNvADc6
fkYFz/YaFADNxOk9QaHLtEQX5BOLGNADSi5qzOgYzVrK+YF9YY8Bh71ZQp+C5FmU/QjG2nF1SWI4
nRyAB+RVId5VxtuNMbxEOIE2MpLWUSnifeGelhP289+bfLRYeE6h9WkHAjlTPFAvSI6XLJCrWXD2
TYAJBatCQcvsqoRdzJRDyMnWl1dc+KtBwXfmlfmYR0nL48vLanS/zrO8VhduqfWFkis/BIqCdgNA
SX0TPuZ20kMQv24gKAc16Nlh/sBaWhuJpClnGkf63svkj+ZK4nu8aqCwtG5CpHdfmSk4eVy88HED
KkJMlkYwg/h2bDUoao1WTFpwAkQFgvhIvFtveyrmaZNGbcFWtDkljEra6L8E/ugboMUA2J1n9xcM
RF1llA4sroOxUCz3pevGSOwro9OGGXr/WsHbI7YsejcgI/C6UZsycis8GlnC0kRzrIBtPTowW2qq
eloWAYD7jj8YWiJ/l5XjagLXhbFQvxWdH7pQB0JkYXcZjusmPZMaGPMaqMZM+BpmqSFM4l/dbr9a
7ePFviZApO24rhavFXXZzIjH+BdcgIte0JB6SKygYrk60gb3w5JLJGuGTyV1IWC2nZSz/akBdu1U
ph7Jo8kvMZe0ARgyHY1sJ9IfjJo3QgRMTSCB2urfSli7y0KWmV9eomDvXdBAWU7stNTjV3Je4r4a
gOtKGxF3FbQvhmU19dNfHCGLVQm7VveyHUK9GkYUXcaQy9pAMsgGQNZPpAOkF+c95N2LoXJYJtT6
QQc9ymP1cCnpA7kWscJufMJpMRJYrPXF7GvDiKAkebSnlIB2sRyXK7b+60SZRX/EgJuP3e6Ge0zz
ssD/zZc0y6knx1c/8LFi5rDpfxjj6jRqN2gsO1UuWDl7TlXkdEIHgwKMcC7yHT3wDwssn1r4CbZx
X/0ntnkLAWFGgOw/4rr9TRQZ86B7+p1uFeX9566CV7ZwLZozzrAua2ARIUceBbzWoQ0ocVroGRUJ
bADP7x1YbP+DtfGfTmINtBKwgpaTP8crUcqs6TIakZDzofcrWuhODu2Stvobr2TQK9/dAqWPCOe0
H0rTQp1blUla/Su/EX1MmFRGlu3QIc3HsyHJ+lj10bZGt+ZHfZxT66VWBtpTAn6iCQdfPC+IIsSP
0sl7zpESr7m2+1xFrC4UZvv+Sqny2r8il4OJy2ZLU5pVGu+UavLG+H2chK8+ojnfXDy6P5pvTjq+
EoIZv3QGse//SO78oUBdLMlIPRuwU7PMqu0qAOKGYM7sDHOJG8pENOTxlvYyVrMF4zUTRu6jyQPZ
ck+Kw0Ont16VODWjKqcmW2fbss7vPB1rzMv345Pj4m+JcoJBC9dMHQUFkLhz8EfBS/r5XSlA/vqu
SVPVOJdrY5N29b+EJDLuRq+k6/Jm+W0Lqd7+AgjIPgAb4ZlNgpibMzJhu3d44N+QhEzId4aMgfBY
SFK4ov8ZxBRFVeKQuz4LGs7Du/yTNQi4+aCZbGrMoQ+veh7HesYirxNQO+brBxDA5xmWQshEk6aY
P+OzQ7vKkSA4U9kjcE60FprCNSFbfrOiC0m6kvfgbq7l8yCh2OchfLbomgomrg5YzRKoJY7tPUeQ
87RiZrmL1rD8NdlR/oUKPtfeCcDMUkUqs33D61IaTieoyA3AnX0EyZC3ihfKfly7erjxO9QJ6p/x
8G7fVP+NSVwnuDk1z5BKLa364UoXH9wdGIRm4+625UWWvFYX1zNk12h0NRzb4QVjEY3eFca2+Wuk
5hBweN/jZZyxDq0H5wFVGdwXJlQOrGxT8HWh4Ov2cjrEU2k9yzXjBKjBP0tDlNjvzRVqNeZKxSjJ
jdBEJwoeHAZCPxRsTc52v7GHaJwo3nPUE8/Y4GhNZbA7URgDlbzvBXjpsVy/CNUi5RfBQwQuO723
DwciJ/ZCslh5LDZIOr2Sf3V6GPp4u1m5UN+ZXca2p8RLUsqADgVxgsA0Gl8esoyu9mbNPDo04/ts
eF8FAjsa+MjvaWgBwgk4TRQrq4SWJFMvp7cXNHIszRHYvo4P1SOtuAKKYBcbwX49o4HVKv/4n0aF
nEqEcdVmkYoqI1xpQgibBWiejZHYHflQNQ+qzsMWINUGRoD17RicpvTbhXr5ZWOlQZDgVxYiDoYP
0zoi58qHR90eSN+5cHE7Ogl91zYxKl80CH36gyCs9k/J5ktVhOi/WplUf3cUiJqBFa3TRuGwTu4Q
ZHpwh+zTXsqPAPAzdKnAiU8RkjcTj9FMvKVbhuQxPir5p/9sjO5kQ5r26NNpED6zwMWruhwCkiTN
N1pdJpzCnA/HCKt6k2qErdFBhC8LZmgPFRT1ZOajKxjWjgPOoRSGZVEnbj1J98jE/Fkn5vLsPJg8
uv727v/0B6c2oGyA7qM79hfX3EpYncQxdN/h03P6UiDxZ8uezxckUf0iBgntYRBMr8ynOW0idCLC
C/xq6aRCtorwhK4jizx6806wS1RUOW6shwllkaHGOpGVnGCPpFPRQu+wGhwAeNJtPf3A8wGT4bGd
9ATxvBEvWHLfnuUSxrhVwOK7LYTIEH8N4/La+9s7yOzhzYTln2apej25WCyoaEqFNamNyeC/ZG4v
sMDEfKN1tUOUsJBnyE+cmru/COvzBOe6/2hnK12m7NlJp+5ZKtMwJ9DpAl4XEh9eOtRnDQk+fHjB
h7iB9HLGwnKUa7RJK5+WdqmXNe6r7+HPIxZufF4hL6FIBVdEbY+Mgwtngzm5T8pdmicT6y8yTfoO
8Fb4WczE7qCFTAeIbZv8Ur/TzNhRha7B4/kob5EXu54DeMhp3YRfiSbJMO7xu2Q7mpWl6p4477ID
gsNEJqERGinYjOdHbA1SOwzRA8ZLkf+5joKN8zsZohanZrHUcTb3T5jrvWv0v0KM1E3qEGQ7rAtI
dlivuOMFYHFbXn+zvfEYzehn6l6nfKbdSmUe/7gbH89KLwqBo9fbrJZ56aN3tleISIdhorcK5cuH
wmaMWocnQCt02K1/Iaffc2q/K8ZBhl5luGfKSflgL7WT8vAcijN6bkDactghzi1XP4eefnbbjYOj
12kxz7B0wTjT2QNA7YOcHwt5Bhv5WuISdlkaat62z2CJww/FnQwsUFAVsYAngy1+JZytKnty1R7e
IyooW2YlCW+gzI6FLtR7Y0+BzRFTDnbARSEmOu4/vcUtnvxRsU9leaNCKz8XqhVEjgwCs240FHL0
OrrStQcCzxLdyXiB4RuZtqf+5NNLLxhFmpSMn1H2dxsXu7CT0W9R14uzjYNI478UiYYRSPDFsEwT
Bgt3Vq6TI3LoyGBoYibX67HARfO+5qOSKYJdo5RFvZoI0Az8rQP1o/cZdsLoELblg6AbBNffZIgT
6gxfL2U/VU8OqEajbM66STu94oW/H0+WXaUzG+Mvgaf3hHy4hxXUN0ePHuv0x66W03VrotcV6EFo
Ax1Wv2UxRSxHO62nVgBW+eDduKviJJIsKpPsKQW41SqkktzIYCGthP4K+0AI22I5roP6iZODGDF2
mHPBxZycxJvKSlnQia8TL8wMHE8mYSkG59X7kWvWuTnSbGqAmGhgkFYnvaCqeaYTBJZpCO82/wmF
YjWd4DmXVrUkhPEvcwNSOS4knct7AsiMGxs8yEjir85A/JrdJnEyc/f/DhEA58iRewH6ZSBLu9BM
t080/29TYUHnh/RI9ti7CMmmJOyGitLuCNX3I/G/IGXA3qTsth2+l3/7Md+BhFO292wu1FedjsqH
0737TpXrwRrGPsIaqgkV1xmSTsFlPAkllhFlxBEZkF7UWJRS1b8uqrbu2GkVq6Oyxx4J7UEvM9l4
R0P6tKFhZUlm31ZZwRBBW/Mf6sAT1oFUsrSdCfwyMpZBc0U0dAnG58gFGCJweA1xGZt2L+C3Fj8e
Mb+hcAx5tzCktD2aH+pDHkvwYB79Y7Bz3GMw2C434iZSuq44VRJ5BHM5YwKAF1lP0cPZLaC+tb0R
3ePiedRtdEqeJwTfjwb+4DDeYe/r8ur5QIxGa2U/4bao4w/vAxT50E+v6jz9TBQ1SNOjj2t/sppy
oDP326OqOJ01hSNABA3LGMBrR1SC/jcA1rWyeVrTErvGcA/KMjyG56ZQC8OueKROg9ogUmHc2RJ/
f2pa2zqpFxid94lnlfnuhtLHOfvSn7vu3iiyFRra9Ygaz83tdZ5GStzLoe7fgUycAYShUiNLHket
FYKRjt5LlMayzVJxa0vhoAvAuZA/0tHXraiZWQciEzCg5Z7M71O1xf9Bw25Zaf9Zd46DpU753FKz
S6ZqULk9japGoThGIfS/HWXguxexuL1ohIbHY8T2QjQNTigDOMcp8FRvgZPivV3L9B5wG79YOreM
a+HNjylDxfpm5dkMZw+7PH06hlExVw1KVcqjXU7XiVphl5UZw9krifJnqT4zc9QPPA+FjKNve78t
0L8zRoTVnQRNCP5GAm0UEhKeG5dUQt2VBS0ooZqg1j0Ts+2JRd/h6fkS3OIJrLgc6ESuB2sva79J
mWSFKxvZEbXAMfyAVX6nLsdiLEjhGzSrzn7R+J54Ae+pKHvaXpKDPwwloHh2tv/Y0ysrRW71Z7y9
IQ8SH3PRqOgjaS2sPkudipSSdSwzJxoJKoUx4clpJWHsNEVd/U72UTof+0KioFswG8VTTaSApDKE
FtLw/KWwKPZBrYL9Ncxm13MLVyPqwYpMBFTN/x8H2+v8wvItHiaXyiDEs2ClIfX07PbuLHA14S3f
rOp/a92MS0ma6RwfUdyYGYLNyIJrxrlA1TS3yrHvVBdtZWQUOfoY9BGJxnDi8MeNca/KauQ8DOMp
bhlZSXa2eCCYqkB9UyWWgYZpcNAr+BtrdTGCULy+qN2anpbyuK/6KzWFGDjpzMiIYlSY2Y3TltY2
DzsgswcOXmPVZ8LIjTfSTGbgRIq8FS/9qxPkYLfaQEXxBh4T5SBTDYQVKCfL7sEAhhYR4Yk9CTYV
fSU7CEVzW0/ZN3rP2SgLEjwZuHJmy9FVRqar/HWSlqRIaKzKl2qQLoMZnNn0U+/LXXKHL69lCw7V
/zTNYwEAx5uyFahE6EDDrmaWOoDNvb4uWW2WAv856KKl01cJTq5XFI/mwjO2JCOan5+9xwX+Whsd
1Iilj4gwrl9knmfWMsQLwxmbkECVSYBVBXAvvoZF9C5NqXUMlsonfHPhdDArojxUIo6uEPJjkH6n
6AcT2hK0ovTRDEl4huISbHmgWIKDmCwELhaJIKH1U67eqr2+bnmB9Y4I2ITTnfWJYbsqLEykN5n3
eAGFrmLjJWBgJzP9SgC4B1MZqx1D74BYs577pbHV54mtrcCD6ySL9VnXBqGFQcXKOFRuwdVJSwXq
s6TSF0tX096PwURky8DGDef17lEVm+PGbspI667HS48eHcloPsJwadi2JoexaqQPmjiVyQT827x5
6nhZzZZWjIHUeViThfGgoVsHmS3o7ynnLDkYWSJlX1hk1f04nuDI/O5D2sVrWMqE5QX2UXVd2LVj
cUddxkslnJj3pQLLdEu6gkG+Oi+3A/niAAYGt+IQCe3EV5/lNuYkOqXwCkInVkrTwFSFdrdnJuGw
gUHCV9mlBBo/yy4oF/Q0fkQQjJEwvOlm7UNuyK7kJc/pSsOnPQihBRUj641/jbwFpr4v6krpsg05
K2TFfYZFCbqnzT0vYHVjp2VnJQYIGx5OKMkZauTsoCgsON+sjwMsboUBqvQF2z3Opxov8NI4wpjz
Vxsti3ZfiOdHncIhFzCvW6plk5L7yIqEeCFNQEQUvQd0NcPxpkLO8m+777UPnNjqVc2GBTynX20E
OXxmSRWf559dD0XDxVSglPCYzj0H+hTC7t1/jTBIG3+fkYc+9HEo0zKXGafwIXuktrOlG+FWoj93
UNF3+tWVM5/Ovxq2Ro/IOZ2+rGGqh4KyVo0hk0yhuRmkPJa9HrbN6A//RS6o44wOaY9bREknZuV/
zOIcUYloCQnqYtL0NIJscUDmDHeMLpOCORFoCxckvEQElQo12uBA8pYBe6oeM7AGeUgMcFMD8Cpr
VFCEssxDvjGAFawEIqTghL8jco2/h/hl2oLmRVsvUEla10AV4+GzT6yOawmZjJf6aKimOf6qdjJ4
NSaKOgZBr8iZzu/XRuCcRi2xfgAIInFtEmtk8LmdGu50m/7OZISIX0pEoETKybj/2DUohUew4jGD
6o/D/UWp/61HRDBzTOfCxzrfRyDFa47ovYoVCht2Fd1zjRAIWkFaGHaXRa9a7xmfiZIacjqtvAWV
OHYIJehGMJr7nWg0IX/W5SMgidwg5pYuULmL9inb3IMd4OsEOY3heWXz3jZXCBUYOHRVyC23hnQT
ai2SNt7Kwlbh+miCnIFV7NXBedIu3cOfHVqDSPMvgOFJAzPNnvOIY3E8WMOmIhydYVHc4p45pBrz
mkHJV/accYYdeEIsjrKnpePe8713ryKaH6G1s2dTMg5VlldXSLsyCkrYRopfp5fionMbuUPXMY3F
Hjyl1t3Rz1J7yZ2st9qdVSpIG+L9ZnOV+4ImmpG6CqMhOinqUq5mHRZtb6yTQA6KQ+zSR7aNExJ2
Wjs7sFK9GpG4E5uC7Gw5GGvoOfNjxwu0STbtf4z2wgIA5U299Wh+EARPTN+1/eNgri9BpXFBoVhg
TtbIx7AIuhr9anZRNnfdsuFsb1n/pbHDOuPQCPoX0VN0XS63DbWZjnRfN0w25wOmcht4x2sUWSQu
5gL+hQcQwMkQ18LrGe17RmyiO56UsuZ0plbF8HaP5fTkcyCakQ9z+sFGec08y7Z6K2Gk3tukHTh3
Ud46R0d8ULpT8bZtHMD5z8g7u0KDu448ZPEBH9oQkU64qyvRHXWR15qlwPFLMMS7OP/AoGjOQqcZ
snEtnQTxnvQGvq7ZMaPfYIZglFwajO/HSV+a15MxEciqAGIfj9wRR7NSek23pVPxgobSvyA54lFx
XaHeJbNTesSguzmhqEU3NjpG3AX3WTdc2XQ6EM6STSB15GjFZJFaGJ5mTbJ3wRITHFCs4MczHIer
fWQA7MhWOEJHWSsFc4ax9kboIImoJ9rL1E5Dccc/VjTK3u8vFRUdQ3WQISloKKiCVuiinyTtQJLB
ggrzcolxW1kfSHy5WfldPm30hryOyKiHUBl/WbOfUDoPUXE8nveMH2UtXZ3K5eGFTPPCvanhuhX1
rjKVDTAKtwMFjSxk5JgKcOPy3vA4CNoQtHp8LsdqEYG5rX5aL3mXlaKV9PdpMGV2SBhRkEG6yNQr
ducCLogDopEPH/obtVsDwd4zWsGhLVnkQJryfVE2zzIOFHQoxyccggYEGFLOKyGZYEPwDDiUzWC1
lZj3FEKeJTS8t8/i4q3D2ysvZM3yu0kd3ndRYmgsbUbj3U5QWxSZLeNOlChw/jTtxmRLBiuG8sss
B2rkWX2aPbEhO3VyhuKagzEnIZ8LksZW3rtOvXKhY3nTWzwFTtitpOxZELqZ4wmuQ63cU0mSF6gw
Zta6ukpky4hjFpNlaUVMFcAuOFMwrht+NrHZVGMeD9yXvh94nWZIjBkfSBIXqfHWPPs0K56Hk5hO
2EJlyxrxikqTn9nsS/lN3Pl6P5iiTvjjzqHsgCmBAtlSJ8azYUG9CxbEVu4t/pxFF3pU79C/QEty
ftjJEgJA5zVjKrb0eCoNyl8dCQy6WyDJYTwDTK5OdfeKN70q+saIVP6DtYE78kiMFkqGrLHL/4gu
woC/ciQZA9OlR9aB098ZiqU29ka3ulOIJIrIDG9IoCaTWFQrRwAxJnzkzCYZYWlH3e1DlzPscDvA
tzHoygV6IJcLn2uxXeFbYYBBZG+iPWCUnCPIOp0nDFaIdSdvyaOm6WmXPOkvHn+9FrUL/6qxgRzi
W04e0xaZGmBOK/L0L8bLiPzG6/kS0cA8YbLrIVfFf7KGu73TdxCamSyOayO1Wl/w9f7F81WI80bA
044nl/gpLZkQgpKlERYuwO1tqh5WPNGL24tIQUaZZbX6ZE0PnptNayYy1lqBjUIuzRl6EIIvnqgj
Ke4cVOGg2/2ygGYB266WxiIGKM823RYfKB9zEZjDt2orBU//f/e087zaSwGqLXEbdekwa6hg03Rv
uh787UMZcgdNrCsr1TEh/NWi2SBJV8+XC3OIPQy7axOM+vc5w4ntomErUulygNJsPuG7gkRE9DtG
xVSJxuXqdozu8mJTLmB267LUxb8OWjhw2+ZuZrKUuS8DRQJeiSlL7ukP0X4aR6hYfR/FPXNdCHXO
+D6VWlmfzxdcTyJZzOlac028FdMv0FTPmEWOCJOg4i93pvyTP9U5hLzPDMq8iXJ6ayRvtlyebF/H
+7lgH0hdDnOygDlkOHco7UKeWAOc1hFfzi73o1bZJxy+jhU5bE/sZAHqnYRVz4ZBf3tBsZgSvr+L
HzVIWRP5GP/xeA6wH0agruNJOPSSU514cv/Qn0UwJxrQ72IqkfE6o2j1NJZhMMMrKEh07C8ZjhXJ
91o/FUZbRhPQUpaSanch0jLpqYlQOdyFHpOQjhHbmloq1MVV98R0v6zNXH5oqEJEkj9E9ID7IwJc
htuhUBhz04U4gShsQAahdrWaiOFQDBFtjEQ1urTvTjOCEdp0DLYjogIBKw8Opcmq+MiRZxfRNLgO
8y+puwqmNNkfNqWfiT4mFt+HqsXN6pptdrjA13VbUat9E1kOWx9oUxS8OAKGSVpsd0NEE6yo71Do
Sb3XwzD4TdmvKenfRB28XUGuwyEaVE8x3cCh6hhbjOyUSPw9Wy8+CUIRIZNX559z1p+MvYA8AK2y
A+TklF8kgCXWA6Cg8DcfkJkAVFwPAdk2qPurIlIP01txPcH1rx/mDXfJfmFQfn3TC3cUVJeXFtx9
I5M6a0e9Yg7S/Xk6+gSXTrQeeshENKMfbG/FI+OUhhFU57hyozWGYYL7gH45168ZWuof+1RfeuGF
UFJPV4NfGkO9HFx4ijEvQ8nmx7noZFTI22S4604iD/xb/ZYo1di5WjSppHXGM2cK8IqJXw7iZsDo
02bLJMEwCa3/RY5MV85d1J5CyoobvktOmvTLiM1xxvlNMV/EUgNX4u2+oXS14uxXOo6r186HxpzB
uB4CB6p3bwgbuLxZHKpzK1a/WwEuclCpJ1HK8RhbRpzmP0XplSWlCc/UuoyWcsBjGbpE6xYbzkdI
4t8tPFHhmDn9NWDRkrYX2lBfN7PbuiF34GX+pv09FTZdTp8ChoPDqRw3j4dGJuNK7e3qPYGHFtBy
5uq5rV7uP8knXty9/Do4rhzJ7Ilm4DPWYqMbAbRU8+MR2gDDGcOBgccb0aNO4Ps+M/XvJMImmslQ
EHBDo7P9+uvA9Kf3fUX8ey/Cw6DcCRA6Lp2P+dELeCLzk7Bh+daks9hfbk0TS2k+a7/b0cdZ/IYJ
ZomxniGXNG4fyDtVfTTSkZ5B3g9LuOl2T8pTnU1IL9yDetLwgkbQHGH1SiGnKaprV8OoVBb4sd63
m15dAF91vW1+Cpi8OXQfARq1dB0Tc0a/ZtlXdpwb1HHsNMR7wwkadpIFFJKnLY87wtRy7JrZysaF
84mfgc0QazsqRO+6ZN/onFwbGDbH1LOGXybrrqLUBXwDZMYXykLTt8hTSC1qLxCk8HDAdiPoxRc3
eB7I8D1Z4t12xPjf18M1ggl1wocPcgH6SruOBH8cITLJDEEknMBJEvsL62iVdNQoreymd/t9JvCt
iSNbWztg0+nZNZ+BeINWOdc/VuXBfdOHRFRcy3YxYSw69I9NrSPnHp8MRLJZH8HDREUzhB7C3R/9
YDByyM38MCBVaONTld9rftLxOJKSibhxSS1EQeuQ6X6xghowqStD7Sv6Y02O4siV/AlOA8KV8+FF
jhOHNRa5MLSq6LNQGZHQS8qxLbV6LxN0unvAkIIwMrMIdUdo9KNVhYrLbU7CoCs8UOFjiCYRmAyj
bRYQCTlSS97pS4xyml5uqt9kvm7HOUN0XVAKs5MeEDBi8txp3Om0MYJ7spDRF3T6iCi3WBU6ZTye
9l/AV/F6Xt/1VDkX6xfzSAaKR3f9jEe5dd0UB2qW35Bhb8j8dLRsPn2IJwsDESPB9S1Xj42OO1Az
zlW1Mb7vJc7JasOYm+ZLSrRarysq6/R0Rto6CGgi2jbPiKNL/I1LdfhP7yTnOAFWPwBONU0buE2x
uWpxaYD2+/CDNjGa+evkMZ7sjSykG3/yPQuE6yjldd1EUtgu60AnGjAqa2ID1nek9co+GVuo/+Yd
xgBtJTmbaMrbQIHdu4+7t7vhAALATUKBTEtPYFpfthvhFSFXURYB+2VUoKg/+JscoHDCJHaFun32
N6kKdTO0L5AuD5c4sA9DHjz1uztksg62Ddm5t6GDjjr0swjc//+XII2rvux/stCCsd8OC7gvOnKx
tmVrTHaIzUq/NP4KHwbrL0XUsGXh1ChNfoi6cRcNEbikjEKGmMMkksx5TbNOWLHXv39FF8BOxkL6
cnrCkQWXTy5V6MSTkYDzxCMEFpNVt/953X2AELNWsD5h4g9kQJ1fqeLE33TXWo9cjtAvxfJChOOP
TyhhxF380w64c96LP+WwVo6CywA4onIEsX9MMkaQJ1tbXk3lgwqrcr9w7dFd8vKdbeyug8lVPJyP
YHd0MWw61YQG6CqRixG9uRVsWdOpNDoNkpTgIBlaQOgH06Rla2VawAP5RbPvqL4TVcC9vy8x0W7u
Xa+BNwISUNxFRZBWwFSIyHlHf/2vpUcIr7HokevRyD1IU+Ha9wCVehhmM1ZCjPUpiRrLeMuDVg6J
SMXIzaq2ivIBLOcv/YZX8n2MkOGZYHmVYA5nnr3nECPRkEKARS3lbocVQJfhWjnql80gX7n59B3R
Pq6tIA4kgglrqoGLVEBKAz5z1Ppv1+WbjcHVSZYBVDuhHRpcgvQ3sPhKN2v3bIr0XKHm8G+RZly7
tAppIYixJ8mGdzgOTrLXeQP3XemnBeKpwZ6NZwNNDHFHB2hM/XycHZYB8LVZzlFLGgIZsZ9AynEy
qruBPVGcALYOSHaCKzw8FGjfpDsyeHTZSk4LjTE/l6d2iRR+edymMfjsLj64kczAT3p2LmiKiat8
NNdzwX54wM/yOhSKxvU6F4Sdr6xwUz/arj7ADTb4plrKvZsxRyuIYp302SgXbf3ntx6r3B8JEU8/
kbQgRyg26i/Alnaa9uzqbupBpl1E6lu8wFCJWxFK2R3tzKVF6q4FUWu9LBgB/UyIQt6VHhkN1eSI
iIKJJKllptJWpj6hp2dKQaB8MJ84bkhwkCAYfGxW94GzHK66Vf8jx2BIvq+g6BQup44EJ32KwH0S
LjS/XGnacbHhSBvNe99/UbbNcyYlGMGYyc8czaYDu4X8HCoUkYdHFTBWQVJC67cZuAkEzr68mAsi
2Cydt/rkpLP2AJTxSaVb5rWmQgqTfIMCqoVnqXaM3qmeyWLqfj5mEDrPLtsY2xhN+BSjkwa+BjyW
bAsXvKAZdDDXPoixbKFtzgkVsDl1r3tbtWJPr9PgBpnK9JNALYxdVC3TbZhYGz3uRW+BSSXlfmEe
uQY+UXnsxy4ME7svpwTsNz+/w+hsjrqSOjoRHEPgzqyTJkyREwHDZnuT+XVxUQOsgNwP85l1IyLK
y1Xy1P8DeUGMGWxqYXE6FtbcFJdNmTAZSJaYSfuAUG+eiYz+ehiD/PwtgB3mX0WOQXLyeoo5Z+Jj
nu6yICO8p3ql2rzhzWPx3T5KME8+2mmkL0M8pf3PkBXoL6PvK+5t0gJ7o9gcJBElHXiTR8CW0RBi
AYLqzVbSy2s8hC9svnZrn2DTBuhEMl3z4o8G/9i9pPqbxT1lVv6KQT9RW1skPxRVPkoOoTgPi+IG
oVW9Oz/Pe5gTGG7sTCePAmibERGVV6eICGGjZzNyNnqODOkE72AcD5a6gnJ0NYtMvKJbBD2gci3X
IKrdRkMb6OlvZ6RIiR3bjF/GaXbxaNTsVRaoxHOwIV+fRpL9RP8/rYGKZcawtTmHy8BvbjwF1pzc
iOBp1TSFZMsRKznzA4WPsbSCXjLnLbXhJaRkdrrslr4FU5rDSUiToew6MkL2PEtHOyR0aN7/k7QN
KTv/YSAVe0Tf0hq6NEe3xWXkeeh8f3Z188Hhmj04XMQvUK+js06lJ3d0q41PqChtvrYa9uveEz8j
obSN3jv0IEy031UCTZwwBxIRBok12UJmgNv7ydLudPKBYXLDYfrCRLvfDoSZkZ/lcVamv8okFnfw
93FtkvYyRTt8YgjhKuHGXTpMcc+XpH7PnO8cgGPWOLNoefIzvHzHzl7sKCiI/emDUaR6HYljodvk
oGuB+8tf//suvIguazvG3eQ1H8GfaNvfwET4jG4EOTC695EhZAVvP8DCzqFNa1yF1j7/ik7wBCjD
2A+AbekAnqT0i4D95luLUyZlcP5KLtfuv/tj/0hNlFWC8PRL72e93ZED6hidaYTYAzOSyunxVuew
HZrr5noMWlj0IwVKNeUcAcYpqPTNhfZBR8jpWMEBgcStjWpWqvLB5mXFicL2Caj3BAjHSz0TqQbr
gnb/85YSJLesB5KoBBvRC9egPCKqwIHHjYDJ93Tn7zRo2Gk4hN2ogFl7YrFnb4Qa88oaQs+MM/fI
q0oC8ptGZc5WacgISLwOTsbJ/Zqz8XobCvTARXI+i6W/WdIeuOAalyiPt0IzUr7aA/Oa+uVe+DpX
ipYtcp1Ft0Ag/Rc2vr/GcsHCBHN+tiFh5rWsnRclh+2znZcFIu2pzOM9d8rS9imXvk3mnyygnRTa
GKpz2Sr1NyFSEnkkim9BKOmSBtN/smpm/wU2uXHjBhHoP2hceqQr0TnV/cOu+h34eYkx/iVTOiRz
qBuMcMCIdqDzJ3jA5ACLVG7Xc58qeMS/4+nouBJKuXPmIHCOAO+1Wvxsyk4OVUMCxR3ZEvs2LqsU
E3M0cYgWNkPqcJYB+WuoUWwSWScQ0JA7pkPow9DX3hkPUGJGdDoLwnve/yinlPr7nYoPmmDP3ZTC
MCfEPmLbYLEd0XkqsaIaAnErcULTIdegnVD90QAic1+7kfCYlmWFQJY5wSiuXLKmyzrQ4suHcxm0
nkhtMTpAiMQtjj6LwXt3+mqwLGOx/iY73A5g+ksJOhTn/zTi7UvANNBD8O2xYnlLbQEFy/+bEElb
XMIMwg/zpR+XV68IKSaOc6kUcP7bLbStInmdLcn3mvC/lYB3kJf7ZR0vHNLVgW3yAWQeAvqvI6EW
RMnWfPe1+Mp3Q466pBFuPsmqXW9RBR7M4WMJpGo2puIO90vBehA+slocw1cthkwnm5ObTNtMEtwx
AYTRflQAh1jJjVEwqrWDtpFS9A2IEtDfNe1gizT6UoBKB5CHRxGpQSOSkc+ZPK1eKzh4yPto8FnD
CiRTD2oUzgpEv+jNt0I1baU0Jt7tCMRHEfNun0Egqr4dBWQ2UdjMKo2G4v99C/hQw/30Ii9tfLg6
EGCwJFHvPqBXrjsRoc6Fnkeh4TPdgWqEpgAzI+VZodSeFwrnPQrU7wgOgyHTPBHIXtVVY4weKl6C
0Qgto6AcglpGw55wXghInpBDJQv52g1U5pNBjm+pJxNTeCT80n5Ga1Nj69eLAXK0UEDCvwKgxWCD
JkixckSCr40RAnebxK8u2n4HBnyyVzLx2oOsaIJswfFcqqkKJqgmYkGC6d+LwyosMijPlL/cl3Ad
04OpVX+M1GTEeMPrymhzUKsjwj6MsNtmyf5D0DuuIUvjC919Skl3cTb/PmIJwDZG+W/dKJKmnm3h
hBsgSk2cjgLaDoLoqOsuPI+sTPM5KcimkJw4rmaES0YBtos6Usjzf/LDufxYtNp9eCLN24GosLg8
szfo9EgNysZcifmUhtuDM7gdUDzAZZiTiB1iBrwncrh8VqI4F/368Qiu3CjELHH8Snpq0PjKqoRU
8dJSvarXz1z9+QqaX0iJDLUsDO8K/GqgjXshaB+O1M0LgA0Y1OlTrBMcC6NByFFzAe0NBnSt1So2
g6LZGF5R56caavHan0ciYjxhH2L39qpjpF/yhqWiMpA2hkvqm8YMiula7D5tkaeRehBXT1Vut7nq
5yrkHhexMDJpfvWLQBzmLMDkxeAyk3YDCybo/cAVIepwabh2FqIwmYUGuQmXjbVMjPnRBCFakw4Z
QFtQ3KUu5CVuuGsewRh/rn/oGXzF8cTjOpf5SZNrnZZbr2Ek48arlWMlNvOAY0RQBZB5Dm3aeMk4
ixEgTQcIMD+37OeZySqyDBoc7UZhrmygCCq0zMQ4CvLwpQDgPgPs1SJQtZcL+WBEsbWTeojI+Thq
uMrMmdMow07tSX5fGsVIcF57ulmHMH0kAfGqRPEpCD3Q5Sj2hrhMySQTraO0iiHX5CgSweVs50VT
h9d7VCp3a55lVv74v6zPeEh0D1luwKd8QsAFV+Dvv5SvVK73jI7/UmVbjXQPClLxWxsqohCFxEgD
Z2Jo0wFGAAmb331FYRJMkIdlKr3tzfQ1MQ9IyLCyCe9G9gumkxWWZLnXvKqKrnVWkq8vlJCU80Q7
a53dC/BQ4em84Dofm7QzfFPhywQFwe0ENdjK/COky+gQDk3zE1UyK/TW70m4Fcj91JmN3VzysVoi
b7xsjudIa53kedh1w3LTYrvb1YbRbIt3M64jj/Z7GuOypBf7XVikNi9JW7zbPUubhrcRqtbgDZ4K
zDCWmidxB0s+qBm+CDhCtX5EtHUZHALT1xbTZe9iv3uxh4Y2P645LwoWvfbexKF8edvoaw7D1Cvd
WrJ2fo76kJ+2i7gBdPX4l/PrAACXIzn8BmwwZqiFohyKLdcBRsjPOKkwsUzBCX+42oV4gdvzwaT9
zstfQEMvYrX6HImIY29kwSlxh3Nb1FIFuiG1+YnLQtXDslvTdO6KQCtOl988EYyYnGSrGdqmrSq7
rxnf5wbDIHwm3KUwstqArpqEyiHG86VU6HEOEOr3Ls4lnxAymAIICRM3ahkuVK1PkGJgtts6BRQM
8yrfOR6YfMBNBjTseVs5cgvHoDZq2gF7gm3MrwsF5xQkb38gp5wi96fGZXlC+BSMDHEj6yb2Rsob
M41ta30huAZrr+oJ2esthtgObW0NBIMSyciK3NjwS4F78RdpFROUiRN9QxbLlkCso3E3jXm8t6p/
afj/0uf0E9L2Xf3UWUjwTi+7jAmLWKUR6pCCDlGcjx8YqGeM/53LqNACbrkPU5IDZzxTPAUM4BaY
jS9XDICIXESJCXGkLSMyxtKnNg6gxt27kNmzVUgMylRLVTO7rAxbWRbdIkM9vuTryAT7ODPJSwL2
ahp9WUO4B+l9rudv1Zhu1Gw3Wqj6RfZh47/yDz5xRKmhV6C/+8U0nkX6wIYBgGfHUfspgO/0ZUWO
rc7vyCB9fjZ4B28jjvAkbzK2uvouqJkKpvR8OBC916Haj63TClYe4FkD0Zy9C4JSDJGJ67Sy0hzt
j4MMjjwsW78+Hd5VxUDai/6is3nTAhMXFeyfzjtWy6iU3/hAin1CQorxIq7rz2kc2X445xBNGrUk
CfM/LrmFPMlUQxhhF6vcKd7Hb1gEMWvjAcOoTv5B47EoreJg48BSU4bvocie9sez0sNWIPQvX3Tn
A8S9qXjQyx6mRaopGvB03DQxZXteS8wx4Wgdj716hDiq42n7ivqLgXAOcEtkvgpB1noKPrU62KzU
tTIWfLh0ARbIc5yAYxhInMyI5feL7bDceRWTRyELHBCR2FIRu9yoa3P2MM+tgN/FMBKNwxxRAlWM
DOkwzgAExBbehaPsxV+v5w95z78PooKofQl8/aSWjcHuN4gk7mIlhHSoOfbCZixjdia/GiCT7hT/
ZVf0m19aqifB+cLENnUoYqpQ4Mii0rImuqeUmCH6SlQHBuqnV00Oma94uqaqtoprFKm7SfcEuj9b
Uwbeo26sS/rZ13V1jOp4xhw4yt2S+y8GPNhYMajyIZaGo+ifqQ/FTG0daq/7q019Sxdo1SSPWFuI
5tWK3CrfrhTgzeJmWdwfopMalhMh5/6HUBliDUfXf7pbjIlvHe9p7ZFJDdhKyyTWwLodjXYKfoKv
LHl43Np+HDrUJ4GOt2uJWrwDsPY4ltThaqowyEBQNKQjs5Kf6MZpkNa5zaE/O1YbNgd+kMQSVE4N
fYakf41nuqOOLBsvn9VtjoseZl/AUeyfiYZ0Q8fqadYo4dw1ncD217LK5DtS8x+voAUUtmBVslt5
Oq2C3p2jIB6JmGAlh63TrJP2qtnfbhGM/TtEzm11u28DDoshYp3gMKQC9YIC4IkRRnZvMvIG0F3Y
T7yn76Lr9Mkmsp5e3yHvLxRESTU17Ijpuh7yozPt/ELCFO4FUVxqX+GocHza1ltkK5iQRsTDoxBA
XtNKH9dnHaAAdTphtsNRDOG4S1IW4Y2Y83BSKvpQ4m8NudBdF+Pdrc+tU/L8O6a6fsGxSLS3RP0b
N39jH32jgeJMHXlKAPS/MAo+btYG6qxFsLav3UXBpdVBhTStlnzBas4nVXIKPdJK/co0CRAm4vof
8qCs3+NvF3lZ+dBLNoQCB4qyU1GmHEo5chQF/9H64izmn7kLlPe+9gsLYUEnkjL3/7RdiawaDwIh
rtMR/JC9W5VUxf2HRwAHKMCEezQPTVuBmiXiLjgzHksGiEr0JaszCp6lovy+skLCO+cFbFX0oPH1
T0N6EThG4EEnvTjcWRSiIrSDz3smKEHaKEGt6aflhwy8SNIogiMqg+BddtDTF5ADmp2ygT4+r1LS
JMSqerPS+v4lXxsfZ2Iu/8LbQc3ef3DaKDRK6M3XUjEWZBCyrSzSrH8hNn04nMLMNUEpFmXy1xaB
UsJrZJubH98C6IGODByWTJOBI3hJ8nxRBm4PEdPlk4e2eYuTrUiuklKXvVcBDk8qw6Jw4lCTMliw
P6uTTm/+N9tt5mwO1Lbi+wtNr9tNkXeg8s8F70NnKIMwt1wtHCcU0u9N3eSLRU3R+A3IgV4FuLkp
Ln8NN42f7tCeCFlcRj5O00hot6I9rX4HxzGs6pyvqGZWntv3FTcPY8B8+GNDvVG+9V8Q0guflXQO
iy4ITc5x75n/mAJlKZ5THq3i0XvhXPTPcgYinFQSWWTcJCvgPUzIRtH68JYgPgnQQOxIey6J+qId
/Uym+4vFzFmT2C1Y4dP8pQ5qO/votDv7W+FfdWYWV21wzOAh/gKwTIJCueLaIW2yQfWt235wCFPJ
lKvChXc8pAY9ajY7SwDsEkVQ/Xf82szvJikNnCPPTD0lCLaodg2LpfACPwSWdfB8JiUJ414dQ8c7
mdmic3XYGJOkT9vTo/7T+H/yotC4oPPSUWzHzVs92WOqNBCKofJASmYlPCRhTg8DkHNcGfPG5NzD
Qc0tS192G8KTFxfpyLBucOgOuNQsht563ZKKv63imDPV0g+8JXkqXCCMtwikXc9iGymAlA1okhT+
2YZVpHsuKm6m1Wp4dOz3sdHyDyNPDesFhNjaKnyV+rYzUZ+19SDvHaHWA80TUZlZRWMES3ZXWBuo
0qfztYc6PRZuCPtjvmfHf8Nua4t7okyxFQ1aafO/56DYMwyvDv+0yWYlaYNnmBZesx505qneCL5E
o/gj8A2+bjx9BknF7ha2YBOd+hf1IrWEGh6ofaTy6SxBwJIocKW7bwOoLIgmncJ2NN5H0zqoPcFr
Wpgp5C/GemWqtYMXjHK2FMJ0Fheq5vgRVBdtPdj3iexue3LdPx4ufwtKzWI3P5ghoczjkKzDBZK4
Nzbm2a1tvucZNRrRObH7ahf2j5UNGOFbjSIjAe78tJhsTbajs1q6EboQW4XW+GvqutPpwlRBf4Qg
j61sby46k+cWJrTu9DNTF38mT58C8qDSxXykGYowbampUvnNzAm5g8Og9V7aEJku3r6GQTgS+u+2
s2233qPrSUZR8yVIzuK1vHjzIouU6L8lof7egCC4mNZS8mQz1iWAWv1JJfkbv7UkHg751s5vZrBd
DPB1SxXwxDyFnQ1KEzZUteLUpQ1++L7yIdJXvIRfrRJaWANSLSux6ybfW6r9tVU3yJ8J/6v297vC
SaGqnISQOLUnybjGWLhAn6pf2eRCl+jOKSSpuHUe8/CMWPEYI4L132iW8kdIcIC3dSpdT3ak9NEt
fF3+gIBvndy3H8u5pFtsF2ABOApnPWeNvBT5H8YSknAulDgQre4fAr2sVvJm0f20DbeDajnHKn5p
5fKiKPPvl9NmxLxPtP6TZXWZkkyqbiZ+A0eTD08qqnzOaOWP2rMbMyg7BlEnNGq/7VQaROA2ecGj
xIwPBqN6v/k9AwCaKncMWSeykQc2eXnV6o1G+UFF3JPLXyui2swdCUFeD/iDNLcvZogKyItAdNFp
Sv1brVd+PEvZNzLLuwoFNDaVxiYai1UIB4YJYjcWQh07glvzUijKY+uCaIgq0Gra3fPzTeiqktDi
K09KjUilyFAfBJDVS2hjCRm+bFixpXIl3B6h9ujwn80OlwWRksXZlR0HLZRKcK9rh/0UUjWyhcOY
lQd+RhMELIAi/McoBCoBTjr+0lpmkLhcYo/2wYBPliN7yOOtEi6BZpFaAnlS6YzC8gf5CnJAavL9
sCPH2bobaaJTcXLEINmotBmL2qNehk+AcLvsoQLqnbLGGy2EcbQin60U0n5bCLWXJZyWgBZjtuqD
Vzll6Nda6W92yM7exdS+/ruen8/IjGfuwHQRUEK1JyDI7HWNWYwkPAiwhsUBnd+X+Qs2ichDyg1M
IbXNYO65wXCKrFfwNeztZPPQ0RZcUIi4Q/nJac9UAMNjSs6kEWRMUeiCwrD/AQwPKkMH3RR1hdzj
l0n/PNgAl7M4h/17WfAy6r/t8C3QpEcZoBrvZGKKp42I/q/H/rl0X+fjwxQj6qjxsKimMdlHqYNh
MmfzadpmljU+oH+AW2eIcjQe9ols2bV8AH0wtfeFBvU8vrjwE1/sTwDlOTa88Rb6AQlvMgslOc4K
Pq24vng/jILspboUDQOd5CWdrLurRwHSVP1LRLiUiXa3443eZk/Tk2igaVDK1ldYdpum4iN8xwid
PyOn8dQ35nc5BkA/iTaugKuIAa7taHBYGZzQlu7lamV0rJg6E0uVdfwnkm2n7wbYpVXYrUR51mx3
CM+ESb5iqgemm3LwGEXPRaYc8J77OzAlk7YGYMpvsPLp8T6ADY71JckB142nYVci11NcKFCZCiX0
BkL86y76XGrsg7sLSoyNCaJxjJPzWzQ7ctxlmF6Qv8bYDFavSbf4NlU+c1oZ2xD6TDGNJF7fSa2T
td/zpsMLuoBmzrw5SNiQcOH7wKx0VMICKlifvDoqvzM/UJull6Td40fbSakCYcSPyemSHXu2dmtY
sflrIDgncc5+1SEr/NtEuRfNqDwIhliEcW4eBLDMnHYncmjYVHcCMfCfhrldY7UolMIVHaZTBv7D
us8Sgx/UinnOiYy078Ged0uqABvI/BAI+2rZ1+v9T92j9V2njpJEX3l+jK4IKLDo0rNNwKLzSRo9
w1moDDubxYQS8gXdbwcd7SxaAhQ5nuRTXUS27nLwYSlHpEUuK8TfxYu2WEcbMUQSy4tFMFb2G5q7
/0MdRDFnHHXIJKkPvQTBKrOimhMRLQHzAOSMIjdjDjYWxaZl+T2+ZUr6L1QaQCOirbdrwUq8rYnm
Pa1CsnBivkky3r8lNfHUCUHZQfEcpW2Rt3pxrsKLDvh3BVfwCuPsPkavowh19k0viovjGfi4teS1
N2Hv/z4VJPGZ3nUsaoLB7zg/Drj3KpHWcED0THpKYeH0ixYGrbfvm5QNRWSNqiiBjSYD7+MfZZGl
KSMs/8eavqU8tg7N1ezQuvMBw2TbbmwEeiKlZFqBu4UaRO+F8h40/V44grxbsqvNu+SJEpoVGHI5
9JFTQvyiPlVOTrRbGVELGnwoZBHO7V8KsoqG3clBdc1Yf5UFEe1WBulOei2BiNK8IzL4BZ7IGCEH
vXCDcPFkG3YPF5nVdNr7isz/vHCe1AiS10aYtp4HkNVIOWSm4rdRAuA0eoTiUbQI3HODZTpLKWMO
cTnNlXVOoam9TvbJfa5MpHWj1qdebygkINPr6teKYbZyrz8bMP0/Gj/DbZQFKP4lVByLu9JaKsaV
WqFidMYqEPf6ZPlVu81/w6S7+3B7yhofU2niY/pTldnHZwqkOPAAYmG6PORH91SCUOUOeHGobw/3
r2ABFivzrvl+Dhe+lj9OlkVgPQUO8MbUc8J40zbaZrbqh7JsIUKUF2vEQUf7AJatd9ELSFxi69i8
f0FLK0gx+QOL7/yNro7sdHW6FPj6NoWO/mmM+2gZTmbzo26DlkleCzddABdGoXg4HiMUvox4WBQ/
zfXBVnKjQx577xatpRqd0Nej9uIHEXhlp+YTNnSRw9AmuNvA/wr0tkc166jxyYNSItp0fZN173qA
QvEsluSMda3AQuHdrIHfP/ujL8MP3kREI/U22txt5cEr95prYW3vYaajhoUynyY/SFXVm8SFOpWr
TWUuN08Pn8zloQ+/Q0SBOXLDLKckhG9CufqIMxi4+XS8hpf6hht8OmTQkCly6zWtyvEk9Gni5aRu
VNUKzpjXikNv4IaQrJ2AZ9bfEZOiPulQBlU6XHCEEU3I3c5In4ulO50cwZVXW6XMwkCdu9e+RBli
hROD+bSAEa8YkL7juWF5Q4mMjd2Go/+gYuD8AwutZDB8d+NvCVBXULlFJB1lq6GbgRGz8gb1VdfI
rbGNidtFTqROM92gdj0O0wtGuTVgCZUe7P0rHkla1NxtgNVlRlN+cd4fmr4uO7OD0rpWeNYcM+HR
W5uvEk90eBv6dlAUTgPknJvUqGDAIs7jxdWrQMOe8WfOWHLv3ft9rl5g81AypX6TyjmAAERLiaqG
qraRo8c6vBkGrusQF/otTSzwNInaV4n/lf7jU0iO4v5gogSqL3j58TFrlGIaj3ZVEob9tFSaUxiJ
PRrllqmsUF9bCkJqiX87ChmXMJqF67PS2hysEJhZBbH4g2Eq5p83hWZTdcuGHI1NOR1xwxyJWoJI
9VL9OHlWREuykHDJFFbfh6gmeKI+6NdJButSr1x8rUMxQ2Vj/rv7gjuV3Y0wtqGvu51iB3KEFf6e
P4j4PUm8zUluSjw1DXAZWL8YhHIwP1Z/seuD1H2vVZjMcXEBtcAjDgZH487uC42Q87aEbD72gFIV
uSAtTKZuF/4hLrNuIgANQ+1vrhoQcEUDbZKwDSqHaC2PQnulr8dwJ7DBzWi9vV2PMj5IDPE9m6E1
LY/e7OPL+KjINuFIdetnLizoPOL++9O158FBHo/AjKtzoa6E3m6P5BC9IProWhrGQ90yvxP478Cw
tTqLJkgiqBdpB5teR6gPWHUQpboZciZD601nzuSzKByhywa7Su3ypAM/uL19jiI3MP/uejnQyBuT
HqjBF1ZP9AMg/JV87B/TLKRWVE7UGOoqVZsWg6B2tMC/zKCtoI6Pn+dPpCPAYkjSZIV8Is994Nv2
5QC6e8yVjaqHhEBZ8/KLxcSSb6hWAc/G5zwxAKEipwWumtQk4ujXhvjmk5KEGjbLgHjtGJVZJcdB
Bxonn4ae+hPhRvrEVixByKt/SsymWgPvCpdcbFgBPAqWDgrJ4YIU61NnrODxFNzhB1U09RlAFNlB
+7zk3g3cd56K6a9Zn2+ErFHfaJ7LNOrstlGl96SRFdmvStJshl4B0STUEO6v4UGnGfEZDjA6FKOx
u7npfuajnZTGIh2EAfT4y/isXLA+gKwgzhRaFv5Ru38pqkT2DZ3OiIg2puxXPyVGhfb1AH+fBp98
lFCNX1yx4eVfUV3+K6NvfMiLQSj8JWZCIYBgW/F0nTbOG//UwW2WtVHVygJXlabAwpY+jp1rz1lT
H7Iw2EGNzoI8oHfcUaEmMZcQzK8oGy86xcvBDATI0jetJgJcMcBhxTbXDFbhPqXaW9+BrXW9mLpj
RaE7HhQg/biWGDESyIAG/iBgwgfqsI2ykQUaEGJk85rbJu8PYeKRE8Nx66dtoiIe+dXYxPInt8nq
xOrCsRWy7WokLftKnUIXQIZ3VrZLqdjpma5QfJeU36eo4IELMFkNlyKS/SFRpXGnWmJcmruoX67d
JwGIRJM8lgsnLTqueJz9TSjyeBW0s5b2XubWpXWv4dKNUOXMPhZ/9cGoYROK5vfgPrd8eOEAlzEX
dlKDwyk6gE5xBt4XdqpJo4Tv8pO9J8+xARB7sFb9il1eu7bp+ufsEgGZOOmm66lp0X3OWdMcTyxI
u7I8ofoVKETnTnKyZ1uSzlCty3sNSPHt8czHA3iExG1rxmG226UhbwW+ZmGyrWFbiHtwY006HNUb
wCewFMn5lU45X88pNLylrNEfEMTMVUrB07Zppz0XDflNXPMhU0BYJuwBCCqo1NBdSDYZQWLWmVym
3hAIT+QBX06xiTgqJZZ3FS1yUD/UjM2K64YnY7VvdMFOE7MRJCXfh8iPpTtpJh6SLvSIH1K0xcIe
vwWAl2v/doDDQnUj4w8jt5Nrl9OnnCjTyDs74jJn21s9X0HaoR53yCr9GhHF75ORsLPU3kVMou0h
mOmQccWWonvgztD6CTs0UlmXAgRIAOPcskxgUrKRNgeeC+OpDrjB+q68tDZQbLgA0WbW1rLHUzwO
1H5aaz1eW6avL4PN2sgwWUvakR2Fr+Oe/oQHrTwh4ODghHKIDUqKqTIHoo9sRoh74mkg5/3XLvAk
TjRiCIhWGriqo6WxcffhU8F+j06N1J+0+rdazq2Oq0mcdkaxCkg4I3yXFRTc3CvH0lDgPj+hK8IU
Bi9j/KZ2OhYPjD+tfwWVuODOcIFtC2N/2Kpw0tsSVaz41RRak6xKTLBy7Lw3FPQ377XzFOG2I4DG
TTK8jVoT3yt4MQMrnp1Pz/8Yzbfw2/1GbY4kXkXLLssYD/NKQjdrXur2nzTmmPWywpZV2Z79v/dc
p/MXs2MUwXGaGWzOZpUrDhUFY8FtC9impqqDpuGbzzfILgTUXma/9E090ruOSGXYqXXBrcs610Tq
2TpdT2irpCf9MVGRsNbgEGkRA90FBraDR1u7l328wmziwJjLtUgfa3mS+nq+WXY2vQxmyFqPxlB0
6RK5lGxgJh6gN4lq3cVqPZ2Us22dRmOMhSK9Kd7eqXHF7OxmVNJ3mNbuAp+FZCxjQfC5pZXOh8IH
XH3Q+CKUOC8GYRwb8uzYKXo0aUyQ4rlSdIOe1FQdScEmnP+PqR16SYhYHgtxHY0JBsXmSJr6KZaB
ANoznseWczvR/ymYio9gDKQICPTyN77jUq5BUB419p/dnrLWOo+pGFFfI1yUeLl3uULREMB1IEfJ
mLaOE8a6oo6Ys7m64qGh0q9Y74icYcDHqloc+0GuRV8J1fL6ynYhl7San9z47cDVqEkv+YdsdlTO
LVle0SmCjJc/wCifTiWi2UPw59sOLufKTPGbIw3pfc1iGJEZ0LmV9hXwOhiWyGsmO8jckSovjB+Z
g9z9xoNysd12eYJ7nj0/uncJL+z+JYV9Fdd5U3mjfNo7GTuXuTDulx28w3fY3+qG0Ztj2i8PG6Cl
hKrp0nnDLQdXC4JVx2W38BVkZYoUZUX1lR0f0xHt9mX1kitTpLilzdKqeAZw7I6a7ViSk/JLl+UY
RJDK+fQ2HrxcaBskD7uRsEj4aEHnnFyA0KomVtZlTfe2IrEBikNTZyHDVPdTwaWz65KYvqGxcHmj
zBXrih8GAathsUgrZGXQWLQXurR1vxdPmrcexCjHAlKJ1birCFxLOiJy6z9qkI8f48RtAO86/sfj
/8to1v2pjEz+7ubKq6AE/H2qBCtrpII0RAmxvzTIKweO19mJZzYElMwYrW8PRUB2wNLcbIr/gq6d
e1Mlrtb5ztmxkN0s3+cKwEuPpUrz6IKAhabr1Mmjp93EMpLiapMrZwKSnCyL9yroqInBULZLP+EI
o/qVrq6TyhbWs91poild0yAmN+oau5Mo9d/UlMlkV5t/89csIHjfI6MuIGsSIeEobbaqsYNkxWqD
GPTZ0NxSm29TI4rpJs38nSOWIgePFzBx1lGOYyKVqLuKTbnrfnkO2Mfat7PXfsVXbT/V1vuDfh7O
CzrrAE7J0Vmx2+Q5AB+ElD6poiY3m/1XZPsbQHUpWPnYRblJAd97o/crIulGphyECTReyeddMcvZ
wodkZXrNMk7Ph2LN52luN3RJUSUp7NaCBPwJpqBdDJVr1iTeQ2nB1+q4Cjt0bBaxIVvEFii6b5Ny
3mSXJFe/15Vp4BLRDZFsVISe7hrRIstId0fpHBPhDIlrDC9WQUSMuUzNO5vEnHh7J1ofy0GKjyoe
dR46Cstl0MtIW3stwNRUi5N0/LQA2WUMZrmL3dfDgKhIS3xg4TetdzYs9aX33U/DwtnUACtoBFrt
LBRX/zHNm0Z1qwht7KBOsu7PlnQZr7Qe7SThQdW9ZFH2Rn/1V67Kqe9EjzwFE589+Man4Zv3UhAQ
9nFA5fRDmvrvxQk9GSqQSC5KVQwTZHpmm59tNYuAxykFXIRZNYw1ss409+0AhRIxPAJa+OvFkx0y
p/ckcBSLnZQdbWefLx8aDpJUg1d02gMxtu8FxwJDGIoXOfKKoLPEh6I4VFsacHFd44q4V1sw6XQf
e3IctG8jTtsdpU5CTUxOuFK2Fyzo/dfFMQT877B2a6EkbF/nYe3vMtxqohVmsDkS/9dMHZxk9rB+
sHAxRNRRcTKxENufAZYYsQ/1BndeBB5DErePwbQY6+nGsYWdSVWqER8GlVJZroCpIOSLqZ+wHzt+
g5qLZxOuwrVCX54uV1SUvZcAYoxn0em/uOWbHgHqs7gJceDuLIJPleNGqFr3kGx41WoVGJ/0p7HK
r0nMgD3QPxlH08LEJfMVJKFcMa8M4oSmSJICkuY6nddzOVyU2IaGO/kU+omLhVazX1oz6SKHUKfm
6B4s7uFt5rMO8WTKSdgc0u6Un4c8Ljd/zOTibd3UpkecdwfhVlNTCAk/5S+FJ/6KVpyRUZiEgdNo
vx8FQg7vMeksDcoXMl20I/saR/y/E6AcpNH4WcVY2x4GrNCf1RqXvRHMSuO0FreZubFrjbNKOg7r
2G8QTaAADwOAyBb0rqw41ItuuPDmWX0O6DQtS3XJJYTBAiq4bGgDaNaFt5Sxz/moygZMzu4YK3l2
2gxvvuyRHuwpJYdxGT6Xp4+wXv+XdkIoXjZT7i8sl1wJHgmkGnFSLqfsctr7R/GCXXi/Ssa3uh9S
oT5HB9zzWc6X8/JK8s2hkmIYMtmTuV44FwcwzaLtjPXOqwr5GR0mK4Lbba9SK9FJTBi6z5Js5tDX
1EwMMbcoyMT2di5rvW7ortZvnYMFrNzW465jNrZZmZEh15MJ3TTwJRlIwfKFGrPJSMBsfOFXttnf
IBHOJdItYMJ+42gdGqf1vZr8X+CPl7FVvMC16DuI99Kfqq4oToNMC6MGRyYXPZ9OiPA18rbZC5uz
rdmCFnsfNRlklmHFNI50SPacdRdqStawEX2f5+3s0NqUmlbJ3+jUoEmZ7ESJFAK4dQcHzQc1W956
x4ZZClkqEPpUgo5GP4HRDMvCWVXMPubo/6p2rB/YKpDgJjjKMVX/4Ko2uOF6XCn+/W/vsz/fNHb0
BfAxH5owWTS/UlPdkGEwBkrkkatlVSVrZvH33CkgBaFVZ6oXi9Z9nZ2VM0CPFq44vxM4cp4RFsbS
D+gD6FpOybAWCLweDYR+F6BuShQ74V9V6xM6KvLXRsbYcMMkzbdVh/6cxvR1hLyekFLvjNf66zea
oA7osQY1iZyfecnOiy/qN7pBoZGOA9za93XbXkqypl7Jkt8Vb3p3G40kWMHFhdRb7Kskvz4g7+s1
3TDUo6FP9mbnpcN2tG/0LCDIgV2+Q+LOdHKSDKsg9h+iKo3NObu7ki7LS7Bh7sjmaDOgmisJT8ym
rIsTogoPYDfOvIiLhciaLVOgoZ9cITJoXlmivVeuN93acMcTWwhDNUJIAUfjomjdtop/JbzTEGVy
m3mWdlRwdKPX8VU/b5GC5HEhNBt8FN3qS2wLPEbOywfLWTZ+N9N4Re72fddO8lO2dzkeCxQg1vKe
d19QigRzQGAbuGbjNwlqRZQ3BpYFoG+g9L/pvZ7GsbZ3Ybu3XKKI3jRDX2dalNj1Wtp0ha/YR1kY
8QmG+sP6Qc2YAIk0Hhtjjn7IYg8uf/qiOpXDDFIZPmVZFjZKVBJXtAIjGf4D8XXqrI1leXqPLBI2
6CSXaFiWkLaecIUuiWMadwKzDYTyfvoh/4CCcNgMVxvP7UR1kVE6sPz/SwU+37o/z2wZJWe9JYq3
cUE/WRqBgowQHVH2HW+VS8Likz2XKz640VGxMfP5/EsSUukpPPmdAirYRVik1OdpblmXGfqBqx6M
s8HLY+QcKvcvSPz/Tr3/sRPYVsmHwXli1gGP1MICayCs+19xjPcIHZqpNJS8uod1ZScdHHQxNeze
v7/YZ/2GKPm1y4G/LDo8uBIkD7u5yTaXT2q0mqTVQxoccQpvRZalrsh0JhoZsgDw0PzBijyVZx7b
XcDR/IndEg4T0oGy2oapjMHmCs5kobUxh2XdCVIeD0YwyjQAa7bzWKwU1FG/ayJjBiExc3ltGnlB
6o/RMliNc8Otb9DLfIvcwesHbS8T4ONyberNiHVIcnmtytzcfIY7TQP+vWIhClqH0/MyMfEPc4uw
uAI1Kk758Q01Zucxjy6UfQ/YeikrXR7TWlkOBRUDS8gJc1LmxG5wDlZfButUHQg7UfFuH3+aw39I
m95su/nxW7uBR+azGOZyzPbgGL8bIAiteVMpfD/ycUcedPygONZoktrhsYDvuJRrJzTldTfvoWl2
A5SSJ4n2Nc+pSQAzksmuqvXZaiHZ8GMkMICkOlRat7wRv5i22Ji6RcFOZFnXF7goPZOdAc6ZyTrT
Y8yU4sbjLBRTh0uP6FjjLwUvqRUFNQa6rYbLHlYgJfhuph36e5klqfNrqJ0qTOAelScrPxA2Ym5r
CogT6EkOuh4ZhSglfGNSMO8QWr15MptOrl03t8Eq4OemG9CUPLNJaCGzYkb4piWewJEPU7KI69WL
xzyAXqFtHSYWE+/flmOyJnnRbx2cpYEWV7q2A8pJ/ci62+AFYEbX0Ccw+Nmy8CVGQZRLQ7Zjyc5S
kH1vM8XJuD+ntFo5ZDXHAIfRQH/FC3NI9IVE1SBUcbQ+37fN/nXaD8CoyGUVCk6ODTV+oK+Nadua
NopZd8IHoffDHKLXUcJiQhbKfPebu5zYjMUkrj2RiGXxBSzWp95Cls6n0NjwfOEIEE2DKYdPW23y
+Is9fdknOghi3cpiokGyqbpEd185I3SHv1F9bbNEtaBVxpSy3RcL59Q7NWuYyCid6xKYmykdXa1G
BjduYbWsHxcYTXyrV2oqQ9M1MSCGosAXhrVTJNFchOAzFoLWlwMauHb1hic0jjfhUlnIb1hPFy+a
R7B76vliCVBmTdnxPuo3aW8lmfSKA71JjYnAenHGeGH56U5FrR3r0eW+Of5zMzOP/Et1PwXyXK0r
gnVa4mB5Vo4bHBXjH2AfLfh/HEaR9T/H6drHe95BR3O1fqxQPhxGyYI1/KOTZOdSlEBH//OHJ0I4
jDBWL69ziP3WsfK8dETZcr1HEI6QDztFAEz4BQyKq/BqtIaYYNDxU0xelZyUeIOttEnwdzHhtZI2
MgknSULUYvn5UTgyJlz2+Ck2YqwAJ5h7zWqXbvJE336fdn3/n25sczputlsamyh/d0cMFXCPvVZK
NbGluQWhFGKyS2UpV5xoAI03Lt+rXOdkasOI0wao7Vh9EzuKCAiE3YvK/ApBLP7mL/Fq+RR5fF2g
S0CjFN5GpaX6JYkOXxRqHOcX4pyBFfWUcrBQLVN0O7xA0S8RYeDhMIWWEAFxzt3dV8zEcd1bHI+7
yGymhm/uk0OPGp5WoMxZLVC0RYS9YzIBDvPcUJWabS+Ox6tYvIPn3Nc21qrbxcJvOgn4cBZZ0FKt
liw0l2nrA77Qfz4LvLW8Zg8NGQH0l+HEDbPndPniW3KZQfY3pXWvacrZFjwCWWEkMJPXMD/VXJ01
8tgy+UuHbUYPgiitw2+LNKiFUwOYfCXE98/sXURWlFCFbc5EX6yCtNyT/nuZJVdgHsU93OJR4/rn
Px6V4Pivl8xPvJXyuguYuMgIu5K9b6Z5waODqZYWCzcLyvGT3OBwz2SD08dBHBVnLAjihMYx/XKZ
O//47R38xkedwz1g5nrkI9HVBLeqRh1Y5QtNvpeNIz2/Jj2dwLOloDsEuCgl7dg0OuiRItAaKYoz
a1ZQBgIkHK3LqRuwk+lopJupXtbXVNbAWAVd/Qu6bSGqv1dWqQvMfz/n74nW0TJwM9DLySBH5R7a
YidICQuhmM7z2ZeVF0xtxA2lF8vnOg7Wn/trudtzWk+ZbP7KyVVHrh4APjTUWFRhvah21am346o7
94AG0a2qQtTIKDaW3m6w6a4K/RzIH547BIzjZQ07HIytjUfAQapCWFHSr5LkZ9pEhFpkQj3A+dsW
eYiE0gBuori1s4bUq3DmM+nsV0n52ll20I6JZ39PjGdWWYhyRK8qg4Vy7sUzPCcsbQxQyb0rvirP
VyspH43l11r72iTV7iL3L/v2OXOvnitdzKVTQuC1lYcAUPRi42S1QegCTUQ6O1XlwR4r46ruyIxi
ud56rwz9OwLJVIxQIfioagx7Cme+ffIrUgSlEE9RFMyz1mW+7yASBzf5fZ4w/i726DbYG8+0oFYd
P2YOTU47SZOblsySj+iQ7hRjQ+WWs7w0rAx4CJfmoVNN7w5yEKVhwv0dmyroiqhTqumjsNyk71nU
rg+oVS21n+m5qVvzvTY10W8HZu7POGh5gExN8lDCydGEddQfpVaE70SFP7R8sEorlzpE3CKRWJ95
KEYLKfTnZadv8rUdV+SwqEXZlhULVC5iTFCxiY4TUA8nKRBVdgWGUegRhs2U2qI19PtpIBONQC4M
PjUn3fwv2yg6a2278gcDQOJBf1u03dc7W46ReDoCRj6ImsQXLl0XWtr0ol8jAoKwiYVA/SOUCJQi
YEplbVh1ddBhXQobX2j0Bn0Mgw/Ntez632jjHMX2cdmQJMXWzxexW6JMCd1d5L2afhvgRkAD0i5f
nlgBFmeR2k39zcsmAtPbOikF8hljGmp7aaScehUu6urKh5f+TfcnDbEjTXPQAjKGjaug7WWgpyJb
sdX0BPiMqYu2ZxRF+3593e07xYoqvMias6jrqBtH2WP5OJH3ZK6hQcpbbLPIJhbRwUa+aGTobbzQ
7JHky6eiLLHq+RRtdEZ+RCZRkJqWqZDCfcLkKlkG9EkfrKUAShX8jiiXJ9JygjVl1MAp22amB5k1
u3gz0XKHXeWKAZz5pJ37ykedVeimnKsnYkvASH0FXnu0lOD+I4IXbUj1fRdM2pPEA+pEr4bBtSG5
pe8UV3IWBHFK26Ays2lboy82mbncvQ1pxQ4GLSinGxSSR92c80xKJ2gOQYxRG7EleHIVdc+GU10+
yXWQh7P5zysr9700UbbjpvFNn3JirMFOfYJ6Db0q6RxQ1OFQvSVLktr9DYeeaDbLhAa/v6/oPBm0
ete7OM7dFzWvCmsK9ZTDwxB8yFesQVKm0v6ounCaX1ZhVvPe8kSPXi2gMeU+eWmr/tXsl915+IxB
eKQFXs4xIvP3MoK5KkkPvHtyxijrpGPZz3xj4/ZhAJNYpNwQ7A1ADOuFpL6tLCtkd67O5/wODPbr
i23fz4cVKm6dQosZyGY6Igw185BXizoEnK3RomIiTh1sHf4FIJA/vCfp2IHrys9f8B0mUWdiRoIC
eQlwEn/NXqW8kIZguyIeE7ct5r/3jcsNOf+Z1teQDblQtf927qUvuRbOLcZuyhYX2+8jyF52PEW3
pRfRKJoxX61uv+FMUxHBQ8P1zSmlqCRRhQ4IDDdysqdk4MVQG0Yvj5Hz7D+pCnx5PyX8DDZBEsJZ
bisHBKbSOuN6xMKDuYlfUKAN8zSlyspSn5FimXcuU+Dux50mr4a31vnv7rqcFHY/MiYDRpHNX/yU
uXHObztQDddx/ZmQHzS9J5yLh3Sa4GngRndkWbFggeJpiHn3bptcd+LWolAk//sclOjTM2ulyyRz
mgeFP3n/5FG4i2sYjoxikJ4Tq5VbU6lvaRaKtzbjyLqOuL9JvItVdKGZD+ZEdbF8NOmJYcmRFwzL
Quqgbr1fVlQUg9/Fx3IaMgvJmKXiFUkTABDJCOqSUMbw5WFoe1IIjXks86B2EFGeCODdTWyussOQ
s0lQ7oGwjKsWnwcQGpRpgnwPy8OA/ccOM8ezCAWb+po00/ThD1V468pHLij97t8oXHcmC7eL1n5v
mEn4BHwgm9VqgBbminryaIVTbjrYQjwLoC2daPszFVKkZuPse6oKn6sy3q5K/dgqGsvn0VIJxhx7
Xa1NszW3tCHBnOBwc9KdeTkO9YnBR47NftyJi+ecVTFw8mp4n4+1S1GJU08Ulc21HHP30mBQJP7k
wAodkgAuG3CXN33MVPYxB6DJQ8xgi4p1WYaZZ/ZN17fG6/PM8mG6zncP8RXL6wLQtrQUpJfZLeWl
Z31DaPSVB0siuFNVrlV0X5V1ArVthaHD/2/1y9Oo2Iu53zQ4nsLvtlAE486au2OrZ+nB3nHOxuRU
kKLKWE02WukouAZMd6uV5DQh+YHsiTxXcKko3JGDh9JCPQ0sH6z4Z7KC3pSwfTUwzlCMOgYAT0uV
rRR9CK06lOblBYwQnHfpOoOy7lnxr7Desuw4fkQ90ARVeDbbT4AMCU5UAkm+lfmnzokjz+BXsijO
o2Tla5EaiHmnwt2k9WAdMK8bTiB4GcLgWZWdgOsQANVtiLF2Js+LemrngxPZ3cCnmMLQDaNmQSp5
043EZBLfKHT6NC388xac8ZlEDyxGBo1lXi53Fx60jvrmJTMe8sYum+JyofYLvXEEpcfNdJPf2nL8
PjXp7AXpgaBcZuOkf1pPPecn28Dd0IhibfLFjJPBcHjDp+z/oWyG6G+Spgtr4I/SAPl1OsYDJpZ6
/Cf7SSji4QiFfvU3FMDwufwelaJNmjI2FivWa8Sswp5/KgCMXZXUPhhHLCCnxZ5EJTMTPIKlFQKH
nm5QlVfMEwOSSZ2MzFlxj7KnqlflfSm8Z8AvHPQGAH9KV1oliRmP1g88Ja9G/uwFxum68tiy5+3K
nHcnqazUGR7zK6tEFziy7WJJ39kkNpIdA6N8EwYXgKn9EbQUaqA/c8wc0VmWvyt2t8XbU/NdXIK/
p/UPjcgG+gZ2XmDZX4XvC8L7G6o8baZlGTtqCfWtsM7+inibAgqYPuC8bh7W3o53CsBX4we/Jr4V
0FTS9Z+yd3ZSq1T2BUrHZfqOFNMAQk+FN49OaQM1uYQmgnT4U56fFxwQ0SSuNmBKXr8hdYVnsjVu
5Qf5wS+ZbgnOwihglPQxnXS7Qh7ZgZ93lZDfXh0vzm5jae/2w9M6+dfHO1Hu08adtAM2acgPuQcQ
b5ArtPwkQab+kb93TkfhBbH9cKkRTDIGAtAykDsWNDZ1ooVqwhF9QUGcCNZ32vGf9HMMRqvhBAlG
AXRh63pvniRDlL9pN4GoACF9RMBoF8p5ssg9HSiA5DDFLrOxOmY76n0ENP0AO8IsZoNFg50+AlVV
IzqRHRVbxF+0tw06/LStTK5igUaPA64LA7aWeAFc0vxPJLrshN5J6FXHkhd7l1s/df15GNjkqjMx
n2428v4SocnFk6ERBSJWUsFb8BiIcsVh7wqtW1xSxxkyDnnGzPRAan4nNZTbzYK26B8NILxzLbyg
b2+jJYWVoYK6fMJTZa93ucHlK9pd3CHxwQK6eeuSoIqMgF6XbKsIO2xTERPZtbyrj6S9PPcoTWgF
IQ53L5/bz1pyO7SdB5HXo5n6DUhRg8AePmHm0MMkf8CyK3W7ei+EM3POOJZvNNuqGXNIt0nkDHO7
N3h3y+6YICJbHcTzjxr7vtzmJkjX3RmDqGzk0Oj0OKCYWUYd1hCr9sWKUSaf1Yr0rW4Rr6m4lZK3
AzpkveXPII6lqyBFqsPbRFpbgahre9W54w3cnixjodEQ9uaaW/TK0CnpEoqjEhwPiBGQO6zrtSLB
tOMu6nbZo3gaLWALApr9v9B05SYggUqlGLkMN/imPR1TSB8HVpim2OB+Pbnv+I8TAGy4Ki7vSzJ1
KEopRfGnauql13y9XH/rtKcJ7L1m+ZdXt/R5XSHH+7Av5oOZUYkoQjLcj4oRt3dbFrKSuQ49EjlM
4+IJPZicNAcSgP9Cb6MsDwRlCVPWBfvpi+3AbezCQ78mO+IiRbHwEvbMiZddQ5gfdMCxyU5PR4gq
S83QCvrnLRTrkaPRtiIVoLJJvkBKbe/YFWxozmVTFHlanbNRj3W3a19RVP2JhMdywG9MX4Nvmq7S
QqYAUQJ6aO++FO8cKkcFHdcYMKCIoSjeoMsbDgOAkBsuhH6ZrkAvvEz64QbddUUDa7OXk66zurSh
aNbNzZMlpyowYs3j6ORy3HyvkCrSNdFwDKmQbr/3AQZp/2wZuogUjcybJYSjBnjvK0uamluLfc52
8KcaOZb01qK5MpkrvrkFjQiHi+NPMPAOqN63P/X5XqwuBxpFhLPMbvNu6G1PwGUaW8gssSw9n+Tq
g/i1qHhSV7YP0lbcrm2oNE1Mx2xdXJ3Qt1iQeC4gW4QV5N8svF3O3BFSmbLhTjoFgR/SDiI8kjtI
b7je6ZSF/DGjtbLJqGm+RR4i764kUhHbboGud2uKy1NCxYz0RKItkiQ0vk6c8mazTVFEyEMwVmgL
B7rT4nnJEVyci1tQB1FvkMYhP8qV3JMbDTs+abYhdpn/6d1BteH7Y9/mhKkNjr+/8JVbeUSiMS4w
RBIhkcZ8xC1mZuiEOzwW/cn6u7UQpzlU77Lo325QC6FCa4Uiq2+ajyevMI87eTp+i/nfZPbI2fsZ
78HyBdyXDEO85/hEHuOLLXNBbGNIkDgPkgJyuMNpw4D4JbhsTTviuw6GIkZJCUi3QA4MIaRVmjE3
YdI86npDh7MKTlhQxGlcsmwjwWojVKr13Dwo6ph21zY59b76jIUYOaCXIptFJL8xVSTQ2pyPnWqj
nzjcu9Vn23yNRw327rzkc0FMsj7pqBdMGO4tL+Zw4IFQZ7fE+ZWOz5Uz0v/b42ZgPXdfYHLz+epH
zlcqKIqqq1qQhFSrf9+aMMGxESH1RJ67gqaRgtSSyTXFluor7+roF8vOq6HDnzTvAxBnJds0FnIk
D4fPp1Og85bG4S617WyqpyH3XE19M8vlvmrNhNUsMFytIk1CVuO/e/pNh6ejVw0ufV2rb/jC835O
a6jMLOD+PJdVTOA3ZRuls8Q64ccBC/p8dbWS210txYjBknLlKQUEMY49H5m/mukXfGyuQkpNhoNl
W32dgTcCymgOvlAhptmxBHDQVMmPR3UJUshgtZWx9RM93oS0r6fCzarG3+elS/YabLO74SCKro9o
AJ3eZvOfcB46hg6DSeDg5bKW2URINctA6mHDEXmhhyVVq0SaYWdhLXdadcqm9nvvsp0QY5I2s+x6
4K370a5bf8xd1f6B+k7LGbcB1FszVftItkpIWsCQlE7Di9QQfH8pQS8GPnbVpaP5n99FhWafc0uC
k/KZFqQBsFeuLVAdN8BE8+TSVLicIs5wuex744GcNQIwx0Rks+FmlHw63VN/hwUf2jFrVuQS0+eT
iQ1xL85IXcN84ahEU8cjLX0bC0ZmpK1lvEH50wufadmYnAvQWAttg7In7eqgoGrqySr96mLAX9yx
D5FCxjHlqzuFq9y2kaJTwuYnuSJx1MX1fo+E5y4mtocp8nTi1Yzzr/ghzxd+lN+sWsaKG3tjcXK2
7vjBDg3wnnRS1U4g1uPgYhEKg2xAFP+/vY7JVwBSdrtMm8yJCliYy/j4z/l/yzhA1X/rpTr8loe/
c/L0apXoJqMulq4UjaNkw/3SqppydtP1X7nyvx52RtBjnoTdVnnuL1uwFZXlJzcDATxzDFOupInj
HgzcGRIWzkVw4+6kxIuKdD1mINEYky5PUqAzHRZLxY8o/qhwzuWF6nX5sGPmvwRiCG9tsYbRZpa8
ntUJunLPJJc0RUB+9WmJ2F6nVZa32x1xvcAMHYFZ5NvNxvqT49vj3e5qY5QPBMe/bE0ogNcW2kHL
Udvw8yEc4nTBAddf/LVhHXxaW4rn93qnmNg1ppl7CUt0Xsrysbd6xKXD9F2qeiuzUwvLhsykRrnu
HHSgvCu1tHIXad5AKeQf2DJL82TRXTrOlxJFmLY/6A1wJsuLHv0L+1HIUYTxphxf6BjNXR50c+tb
8AfOXNfQjl7emN8nrO7cL4uCQYqDOvKAMZRxW22pvqR9OakphpDAvBUwPHboZVapzNScPnOhLAuu
avnr3FfYVbfefYw6YbR6HUMef2WuFoKb7uiXUgnIfD7eRC6N8eqjC2cJMIVyCNG9YmfQLJO5jl4l
9g0FJEPAmriLyyZSqz2YDA9djwxLSNh9OVZIRZ/J4l2r2fNRLfWvQ6nQiLiN/Lnrm8beoJ2X6djN
yVEl7+qlbY9KgfXE7OJI+EkIg4KFKFMkAXzzloSSvvZ1FQB2cwSCfMKY7rRy4KXm1muxb9yaNqup
WuDQYR7l73nUxHqkeCcWR2Dbon6HsIVmIdIyk5Vgki6D8z1plUXjszCiv4c7OxTNgF5MVRY1jGuq
uCeSCHEi225F1q2Ykivp5oF4SmAvj/P2SYYrCXb+Ta+nru+IqwajGp1RB5NYY/Nmxd67wen2laNo
fRNJ/Kn1viP4wUvyUv39ELCXj3lfDRs6KmBBR/K1s9SZq+cGN5cf2TlQFJ1F9pPBveVsFWWd5989
Foj4m4s5rQ8Sm14IsGqje7RiZUhwS55TV8er41AtTYxXaQ8IIqjhG9QETWUQmNMlDOeivMe0cCUs
HByYJrZjt5PjDneVz0on4ltbpwtWDwCNCGqC6lcwi1gEoKzYZBmE/X0yDGRFfu80/VqSoxsXW6Co
ZCV87uFNLQ/MGT6EK4uE9eHZf3Ne6hl5I82r1DVnTL4A+iaYvwpa//QTqLwgxNmdkohi+SkXyOXH
tDD0CP4bW5VOAhihQP6uzJwAOWESAGSAcWz/JvYJbX4NCW28bM9LfJ4bzbbwjSew1+8Rwo+h1TB7
yeeEmIw20h+lVYhe+aU6o21hjOIQm1XO9Jj6KobYKcQwzxrrm0l4JuRb9JnNntpQ1pTUafPYPcCy
8tRjc6tpraVd6zAYo2LGXZTxVKz65dNIdBCjYtO1z+nBvHOSixfekucWtKT2fpe8HmiicsXF6E9F
b2fVS5VKRmCEycnwx3ANorWXQKPuIOxIQBDRaDV3RpJo2bwg7vGoSZqH+CaXsjxgWFDzhqh5snMF
KFyavoA55qKx+ojbnuD9z1gIRbxtpf5Hhk1qfKIpcSQJR7cyeyYIJMg4hQE+KMg4pl065ukOKZoO
StNuW9K4/g3wrYmFgOZeK/lhXSoVqSXrz9E1vaqJ8C784n0d8g7Wi3441TFtBGLM4Y1acncXpdhP
aZg5HHxIifVukhvHJTDArxpVGJsPwzlHv3x8M0E7cXlD4CUvTMd6d7H9SRg2MWLDOpoF0wiBo3KE
41DpNdNmnFHWNB4XceKI5A30oElznK9FHS507q9SUkBlZ++DwC2zzqSaAMstF7M0fuduJUvcEYzs
SFnn7ABEtdnkgd45BBXgTfbvHf0Gys84Tfl+6F3kPWv2JzMUF4WrFkv5bOR/22IHgf7hizj8PIGx
IYU+1VASNE8Q9celmzrKV8L8Wuh7nWrSu136Beu2wbyQPbFbVm2+CGqjvSupPSUT74a5qTq/5C0+
QXLpOxzeGayhX0wybnoonGWh/6VOtydqQEKmPQSWDz447s6Q7cEBi1YvsVr/K0kLnD8JqoLFhuct
IzcRgEU/PUJGuzMGslYJZv7ArB/QyPBFUD8r+DBbq1vZ5MF0xGkcR2dc+VwJ1cCeO05AKZ9+s0mw
KT1aI7aBLLwxmSmHFlFaWgjUaG6WhmDvBKJYPsK094fNY6nm9lddJHYYfoBCzOqTZ1TYb6ryI8d2
684JI/qodp2AGvm6U/7e7dQEuNvTcFErJKSYrBPk9+MRo4uBpfkqhXe7fJMuZ2pxL4N6tLiy+tZi
56nEJqLE98SlNcvJyUraSFPoZ3j+hmXaVsNrLmGXw8/P1fVDpMWKa5Mo3PykLewIUnHItbnqL3JO
uiAEg9MNWLumqtoydIvmrHhEpHzP4QyDHaPPxS23rmM/1hqUvl8MTchOFTlsldHjinP8gkx1+HJL
/lDY+7A7rpsgIwfBm7YlpKMhjtLwfc8BacAtwcgHypxdhugbJYjfIm0fxdP28lvdokWZ6iVO2Pag
rZHM16aZN+2W6Kw/KCQhmrzK88VKS83NzpHmIwgiYYyrxn/xGOicoZBJs9ZS86gWYYXzIlvnSP09
xZFllgn2oiTJG/Le7R35XQE8mAqZckNeZ9koyL1tGdDrnHwAMaKjmSlI8mD7e26WDA7czjQUuEd1
ZVGRXxTozpnXcdIuJLUammEddbd2IKe5UqaHHzDKP65xaXjcxpmGD4wneSV03yNPIvSqLmctXF6z
WLV897Nt2eMlAUAO0iLQbGiQwzy87vyfTBS7ATnVW/hH8Rg8OaGk/s8uE7tqw93UWF9nFWMOj64A
Cu8jJomBTDxSdV0kbnl+v0juJ9SvDUQoVw6/Obai2lbhTeNT9ELxL8ngbb2yJUZVzBpoDU4LUxd0
tf3Nwmm2BCdYIlqopH6HftQk7ZIjnLkLKBC3WQoRWfffCCWRV8pwlGMRjxC+XE3S2K2iSJf1N5zM
xaw80JYXYIGG/o+Id7FhjAqO/whqhYrtnDVKbvKwOiADFzzf/wpfcjkhGaMpwJYSTCFr9PTx64Ai
OAvFlz8AyAhZPE/TvpUQj/HrzIMKmaI2a7KkKV83lLbtu98kBDpTT3pwgw75R0PxAWOMYowModas
A9gLcMGbQfZ/qbq1GZmams1SaAJdF7w+qNJUmdvW6PCA+SKhW0iVS+IQSa3toe2Xi3Fl+67sL8d8
gR34rTtZJtTOovm7FE/TVyxa0F6hPXov3RYCmQWG7cn742AuOKjWShMlgUE8OLReQ53ioDm9J+P9
lxHljMMUV0QOOiQsrWp83g87LUmdoZaw2NYrzI5bRSNKQ5RcU3Vwi8QyUUamw1Xy34dp7fwNZO52
1gBUYihy9M+Ucih2nUg3pbl+TzCjrRl6P2J6rOesbg7Gac8RnbhWIdYjoI4ygeH/iexHV0gGWkf2
1zPZi3fPzh4tRc0PTA+qKx24dGYp5qrWfakDAvj5vySg53J4fb23LUfi+j6MHiJgJAU5BtCC53J8
fe+U65ksMCTw7PG0BN65ppwjvMp4kLJwxsI/7c6pS60ZQ5BbNF79sRb8EzknYqQWXuTnKNtr9Mrn
xMxyO6U+o0RA06s/Y5LTxHz6WUKlbtAE8uK/CQByL/hmcEUuLVUUyfwZ3OYtGnCK5/SPhicrVg1J
/jf+/06KGxWuu+Rm3m2rMpGhZD29oqrKkJA8hdE3sq7LlVjbrX9qOBBsbN0ktwMGnB7BGbEkDxPk
0W9DQLd+0fa0ECmrF6jvV/DDoo17+anZ+TT1PeqPvjsfTI4PfXuKzqDjfrtuVlQZwX5cMDqhH0rQ
Dmlav8lDa62+V/Ha2EEQft5xX7CPYEonC8NvFtDDU9/nQzU79hTUEUWhAshC/EewxPhga6jD3p2b
J2pAe0ezjh9v3tprZ7arON/FnxamwDoDd9pmPzhHmecvVwSZ9hGBwHxXtee+qs/gSI5bI4VD1WuY
ejW+BPWAVMKATU8QLstwdu+QW3il55K9UdXOeQ4SHA0+b/PzNT5dBXNcBkhlrUEYkzWhJCd7ye9F
6JyW1wuR7/IWtxjFYBivPdF7rk7tx30LsZ85il02H7IKFZcvMt2eLPsHW2vDlN6k+3Dx/iMmJ9p7
6uT6ssYej/lQyxDq6jsRAk9cZ2okqqHSpci4wOGc2cUXs0Q3AdqVxv6tYjwcviKbQt1GUoipeazN
6sUTyVLalsjBreDTwbPJJbOFazWMOJYVjKMjPy97BAJxfIp3/kIMk38joma8ORqe+0aqGb/1neoj
dPyDhTAHqgq8eppkv4b1iCGvyUwkhjXNJ9GZ746I/Uw6thscFPOu/7BlatPcJPyJr+g1rpUfwuLw
ij3IVxfeNcf5MvNCqJZ3kDkHzc9G8212LVb70ZdrYJLPc5XUMbpR6gvdRk0dKDvHPTp3CeBdLy1S
4spQc629wkuDM80f1EhfcjmscFZZ0Te6VRpzV8/8aXnm0TgPh0zYrYvEAaWf6R1/ghvwy2A8rOHS
3isfaRVOwP3DmYtyOg4mFdRWxDfB/Hf+H7RqW3tMgg6mlJ1vVA01AEzHFUdQe5R4BK3U/5+qoTTv
f3a8vw9qyRGwEi93jWLmdY7oYYRHVZadjoWYxzhwcLrAJ3ui8Mmzu+j0vUNKRfP60Yxe60JkpnmT
hauhEzFoAFq1GKRMiWrcHFZoZNE6ygJv4NWsChgsknxNBGrMrYj1FYedJrnAmSGtIYwvL9g6aDqW
iQ7jAF1PxCshAAKP+UCo9yQX7luKazQj1hMNabkurS9DVrfv61jyK9DeZbKhqVUwa8tgIFciQnC7
SP1tZ41tCXS1paosf9960xxHy1LI3FDMpDZjfoW+RGEfxxmjNhiwfyAm0ZU/Pact1/r7PxhUr0x+
bHij/WZL8KKK3lJXJGppMEi6d2a7//yCsGWZrHVTKucBo5wS42E+cRtuBzQAgJuHVUEz2OLsua/W
3uzadRs/pZI4GVjWvY+GJ3FVlwl15WhRQOdTTb2CPsT3Q+/IUsspcgO4dgG0ig2e9mQeR0gtJdpb
1zHg5IWfpnq74y16DYNmAcdNZ4h3g9XTlsozwbJ/dJrRe/xDiEOGBswlM2opyOYCJtklmivZ30oi
VEPpnAsvqgDDYHficXsdKY4XTaITpDGe1j7kekynAbiek4mAdPqmaiqBLbu0dq7iADOaqDgnM8QN
5riI4toiGB9nk8/O3IO+xKkvVm6og8RixJnA+FwknDbD3Tz9CKXMo/L3P1Nzpw68Nd6GHypMyNEa
SJ/bw1Nhnpu3jfc8Fdi05EcgMrpywkYN9RbUeUqqbvw7Poo1wQy8mxdRQa847wfb3/qgCC1fdRbJ
cR68qjWXWPIIguB3wA9vugA1F7Jcs0Mq7bhxI7mXtew7YROQ+eFAd6XYYx6ffCZrWWnEpBPpc5lO
RQCXWrSsOWCtkA0B/TtAUute0yapsgDs3+Z8ITrA7NYY0XFZic5Q3crea/Hi4BkepYY0myY5Zj3w
k8eeiajP7LcNmhoVbEViGKsKGMbJ3iaoEfhqqQuRdwQw2H7nKd/lcMSCVAsDviX1o6PN9hsG4WOr
9r2+CWmik1iLOvRDabaAA/BCSjrKDDZdOI2dUNCstLNv9bxX3TqQYP8PYGk3j8O3LW0cfSmQhkYK
JyrgxWVMCSk8WsL1zFspdW2tNV3yUK/O/zLlMuyU7X2g+JkocWpa9UZjfwlQIcCCSxgj1FHgpmvO
EBMcmy4IBqmy0wpeX+Igtwk8pZCAUQwGnDEdzrv/jhS/dvRpgRZSIvuonmXyIbPXSDze+M/cwOiU
fXbwrn+f75tKQD28xnSnS9/HIYa9vM2s1kPqrqREX3YltyVqz0rGnh1BunvW+Dx+Bj98R2NrvZ35
okolX6JHvr45NxQf6O+uLeO2Y09DOA/MnDCFLd0DMDGuOZyaK8jZK/1KvCbWDXeQYRp4i6unHYh4
9Vb/1jVETwZuxs+pOdoL1HI0xk8Qo1BnaBo1cf4DsTaD6jt8XkycXNNQ6mFh6PA9aTnVon4rRQkT
6YhT2MgdvurHv4W3FhUTnoVN/o6z3OBiVUsR7I+TjaCKBn1QQBRU7h7i2mna78CWWiHzussRSGTd
uoriuVVOJQrLmJkaEcI8EVfla/mp4Oe2l2c1WHTBjCEvCc2i+NfPhmNUEtRtCNzYS8WIH+lf/Boz
Zy1JYiQqpXtfAsbojGWBqYiTsvRpngbbWdkpfB6oAVEcPOKCHnMteAIUfgUpilj2mFYzEqiIBgfR
H7wNNSQlrJXr7YXJdaycwlVZQ9H+r2ebxZa+E/BBRH3iOBMERpxvEFf9r0OaDks+xTFRq8W/l6TW
liTpifJ3y7WcKzGHyFKEoPTrudUvtj75ph3POdzjX4ETVK8mVJB8suFPIB2KJYNEHScPVlkrrpDm
JIN2DLAnlrLOyp+157AmdH4T6q4CLU5a+0O5xMIniBcEgYZO6pOZbt+2yG2yhu7a1xrCQckiqYjp
HIUw41prEHPDDJRi1Bj2mQkA1kicCEi3Js3jMlMjKGx0ZJVPWi2c4Cnd+yn68hkjeutjgsgd3tNL
y9PwaEEuBMyEzlLv4wyGGrOXcVMYW6rt0eUwe52Kd1ovoXmjNjFrFu5jr/QfmeGZEJhhqB8JuV/v
NOQwX0h8VRQfs6jq3ARrlXPMlw+CY82Cq9EugeamxxnblQkVX+BacJti+zov7YX7ZyvuaV1hY68k
FQfJi8qTPth/zYB7iH+bxYONn6/OemCvBf+Oyv42YZfyWGqpoesH0I5XXKgZISx03U/yghBYbwVR
rwd5B2LIDOVuN2IHVhBb3A5zqD4Uv74X7HzolqVOFBDdqnuZc+Y5IRg2ll/YveiB1rc27u5DYgTQ
ilH5U743h0d0RUp8ykFXjqfy/dig4fkyXxjJcTzfHngkpORi1m1BR3B8VaZ4xIfjU7hEefIZ1e5z
CGeKNaqcfwKEgsoDAGzwyS6GWAq4SO+twjONBnwFhjYgDmWIE+m3eokiJNjC1W3v/lSEzPT8SSGU
R7AdwvreGVUJYu8RXojKmP0aPhVOrcB0vBwbNCRnIWT4MXUMWXvQYUbfHpewdngfUmUhvTy7FJyd
H7Jbc0wbaZOPH3sgRtm8EkLiXqzRQmX3Z/5co2QJ7yeRWhYG5o+7hZJ4QEUlzfqrgkfHcnMePLJg
JnnGwlJgckyMoLFA75eMpc4raCr4fmE0737XjwitaYE5xBAoibK1a+O3Wnl7z4nniwkocr4k+4P8
D7tR7i6XImgGnPdNsOfPZUR97x3EyHF5NBg8H7J3RZpdzRhD8JdCNLW6WN8FRpIO6h716gcrdvF2
2xFfCMRSuPzpzM0nJHp1pCAT+YwJaUZZ09/zcnuG6KdSu79vPeQEPDUjwAguh3h8P09UVUWZcEcC
Fo/4M5s6fj+ADR8xSu6fbFSvNxht1lNVykadR7NW2JaBWYhwZB75ZK9j3D7ujcfeMo+LJjz4TcEd
r0C7dpzdhqI1tAB06iYHRNmPAK+vizmA1wHJgoNiTS7DBhGmxNq9EXD+IVkZm1akDVJjSKG49nIu
5qcOCTh+ysm5VBW39pLQI2osOvAYmG2GXBCM11Yf6d54bjhSU78sTnfkl47OIzAq3CJlGBeIraCc
0y0nt8IVajANnNV0a2Re8/kpZmlM76sp6+WBgzTdpIsF44UYGzcMnvMnS7lf3dr1dLurUtL7EUc5
JRhKHslN67am8W/euPF7N2HfCznlY4QK51pxPWTWbBeHt03Rl/y9F2x5eU+Xh7QjZ4pouPu8Tql6
ikBCNx+h6DOHpUKL0CL7T99Y9XJoabprIJLlng1MhTbTwT/kxMnmTO8KBTB2l4/fwPvw0EYfttjq
2h8U+DAR26vmBaG73V243XEBQosWyP5qU7piOuVBzkjcRAKqoxb9xhpPO6NH40J0JTFRmdO7c82D
mm5i34useP+y8JXoUpJcLYixeF7xwDHR99Va8LQZfoAQCwcfjVW6gMaYb6f6WkmzwvJHEIIVyzIt
pgTwl8HEu0ikNa/FezbcEeW3+eyh8ih8Qpv1MvXHaC9cBdSuNtZLtfras6puDhkNCv6Pf2Vujdi3
chrwU578mMO0pBY9YZEGwgDmSGyLCSnWIytCfzrx1V4WENSPNHTMYnJJk2T1UDbgPrBWbZn81ey/
DXIVeCr4cF6oXmTvN17gmqAFMWWPDBcy79GJIHyPNR8nnHNeVfbNzmMCwm5ddaTaVWa+NPd2xTMo
uom9oQ2h1/XEc+A53V4qq6HHWjmfltWMQ0iB4SRmytZld/LqcJ9Tkv600wk8vXxZDCiG6SUnOWva
QWu3LChuv1mylWPk7NOAGIsnqEQzzWuoogiEDl+hH08iGsdiWdpXpomjI2jHToThufVu7U00oYbV
8uEMcVVgy4DEU4aAeK5PZCci7kUg0iZ2vUNOqKKLVbfOrq9zBBoJ8XNvgut3No3qbtPhQvcFMiZT
3PwkaVWyBLAZuRVnfRS6JuegzJbwRtj4s/Mhf9WXO8jQgiGRU3rjSCcJTuG6q+wyRFeCSgYFVy0a
+fvwIa1+NlGR/W8p2+o0jGBD2Yj204TRYhLPobJnA6jffz5VYYPMIXCkCEioz9gwBmuMf4UXmEpQ
7THd313bid12GCNDfReadCyuD5nmIvA2+yNm5HeLYmQnNEWfF9n1q6QBTGwHvN4Hr2Ghu7zb+h95
eNEwUFXB3IMxK8WrcG3bxKb6HR4oeszh9x452EShZriWCbMIXdYoKbQc43chS2c9ojVR5KGH6zDn
8hEnhXfk/QrfMW0uc4Q4HWhwNy/oVe6RI9laD0+LcVGD0LPibNgx7zoU27q/NLF1SrEmtuKzjP3r
oN4t8I2HKRbNPiptOz7cKLAiyekPiyjz5xxxoYT28cOsKo0vroYtJ0kRw8H2KngCJ2QQFH75BE+Y
W9F2vNg+OCQBDh2btajYe+ENCyxLIRfAmRcEstWWiM0gQjDWVqcyF7IJEKogBWT9OwlgwrvoJcgq
wM+DSkzYZxVhothB4FW0cazuwRhV1oddtz8wyIiLC9/GvOsir91H8hMMwrGs/8NsfNY+7av1txWt
JDkHzYUNahkPPEUdEZqR8VnbM/DXbyoUttvxJFbkVRlFk4PAyiAnZHJdfp6yonO+RN+u9KEigJts
G14GhgH+FPbQsuiaJwSNrkS6l1QbVSddKmMDnnj//sIVI2q0xLWIgC5lI1zlHc8GaMFIsewfwief
wFluGgZpNIuE/nR/jJQ1nr2FflUja2sOnEwnvI7mQhBAVL75UMY5WQSDr0C5MuGkYMycdaQzXqrA
F6YqH8wFuxw4hifmwOjA497j2ZGPSlCtk7i2f3J/EKIF64NUnxVSZZq1cZy+0z3A2/jcDzlDG1Fd
gt7lYbP2CYwaYf/IDqp5SleMBPGjSFA/PcEYOm6N+fqrDh+fZgdWcefYYJVwH20lz10fCwjrsOfG
dE8ZyAKXZdjSUBQKlh5sjbBvX4O7mXj5e6fHHFpCniKQTTeHS7ZMTBhVS+nD6CWVOi1Z87FSTQQe
2qKdlvXJTxbB9RLFlEXG1w2JtGI8vxlyCfA4oeMp9F30aQFW5bRyo+Trthm3Eh/AvcPWXI6R+RwQ
X981A3dJtGp/2ADwj7Sbd1om4kTFB/dhvxbIk8LSzya8hoMVyXepKrugVnqBQ3iOBo7J+dni4t7e
17lpupEKHFvBH+1oGExYBsM6onvsKiha//Wqdh7aacDQJkmY0fE/QxGY1lK06WWf8BRf6GHNJBHq
SLei5c+6r3tx1Sx43z4ixDnPevEES8uRQ6JmzT9uPmbDFrqMlWkV66XaYyohB05qZlgIOMd0snZg
ONUAv3cGdeNMl7kEJeFToKo9Aq1GNprCHpkVxoc4lTHuSgJb4lE7XCNlbyDIdypdlJYQ8XLMF5u5
L6yEYMRTWqXqjPYoaiKJvkHdEvMYyYuSCxnWbSZr9dF8vP/7HQpwefxLQ4pLwR0HGOgzZmJFLwUH
GewAImFQV4ykNC+kohFAQwJegLL9VbyEIikllVCK/eFNFADPdLscQFrS7S8hp6KFxZCrPuTvx8op
iLOSire1dFAev84BLBUCxc4SHZUP9ADX8pUhSPPFwQti7TUJRVQFgss5GbYlCNYUDmxUsBobZ8c1
UfYrLJx7ceRwTffUxXAb+wVfj+y0CatSHUatXSmaTaHOHZ7JKZP23uml9Vk8Lu/W7q6pG+0bzaGY
cXFWRobOCCW4bwMh8kWsDDE50fd0H9IaIdDXS/GzXfE31BqbWbAmvXpjfTmPyryHCZbBXsOGp0is
F2ZXeu9swyGl8gKUC2JSRn9U2wwMgzD5cBWo3eSM7OelnPPejjU1wAJbqzdZAC44rExMAdOdbeME
kgsEIo9fFdrtuu7P65R2HbetMIN1baDVilXk53n4juoVSm2ZVA6FFtVEusvTQ43rv04+mHdYfWrW
LEf8MRMzR7+osDKNnO02sb6u4gAEjuv445sw6LwbemX7VtXJjQzgR+r+iZDzla7LfJy4t8ljBv7X
ER6/5/zA2/N+bSG3r8YIr/zq5lNVeCabbYfl9//xf2n/YzfCoE097Q5xzXNWTjMnJPsBPiTdSMvo
Bq6hHG2/6SckCVc3rRtu7ExKIKr+Q0L8VAZlTopw1mvfzuEMB/ccTC2Eo7XvEtr5gI5z0KamY/HD
UzWXgNXyYkQnNR94Qmq5K9Dz+L4aDSi1a+iZyw7kj8HMcO7IipkIZIjMdzD0zL2IsD23Q/juz3Ob
XLtb8/+Gk8rJUv6BMGoP5ptoK9jdguBmp9ewNaioEX12viwrSV8SJ9yk0tX3GE+F94F0PurxXzrG
sFKk0fsuVlU6wLGh6W/2qfbVxCBipJQmcQtDMa2K0YgtlvygVHD8oZ6A+h+KyYaI14HfwppiT+xr
PaxXjmcMg/Jw1FoMSdk8s6AO6SsqEzg+haKKfNdKqDWk6UcaNz2RnQF6z6S2tNl+qijdNwvKZwYK
IOnLwEAgb1UqfQtUkS28Hmvcp8SF6+ckPVcVp9XEExW2IBp1RE5yc3BQBgZNS+JZkrHZPFf82KkV
XiDqG+n5jLR3RvY/Anj/LSuHdQOfa75rA0FMcPxJ6dYM0SITaNDI7UfvRJ3momYl8CX14ee02z2c
ehvPxNhqVsIhsNp+S2z1Af7V5OLkQyu5cODy99dtJAb2knVBj3vbDI0Fqc+0OsU9BHQAGQ9QTA3u
j2EfgBRokQfk0QXD/QiWD713EiqbbvZHTUVHfUFhOVdCux4+rqZLUPKsDBV+73GG5XaGtvwMe+uf
OG77FGOeaNw45pGi7QoME82BljWmUlAgpCO0cRnQChPir9VX7oiUpIq+Zn/HqvRDCQ5Ld9uDeDg9
orh64iewVlfizj3Q+5joOhq8Eq5lTfwafadJlmekNU9Ov8Fezq1GLEGgYQmXxBV1I7UPy2/BuZZ1
2O40hzo24lsDCHuS2AmzbcEWPoL9Z9c5mfU+ajQeQG5Y/c8oIQbRBw+t+/lyWic1jDKy5QMNCske
vTIZh6av/C7koV8q0mJ5QG+BcI2wiKS/LUFZftLyt1y2nAKqYDPEhdbrqMH+ySMk4Bf1+FP180i7
li/k65O3dL8OnJCfNytEJ/Vb+UOCoJbwqpsMukczrCH5sOZuT8yjzzcTcLGc6N6/01+N4P/2geWz
p4dD7JS/7vkjcuw2XMsFkEOo/OD4OyMGiEpyTcgF06LtfCbMbHX6kXXh8imjAxmHWl8k4F+hP85s
i7m7LKz+okGpJQ45HJKC0Fgr9kQc20RIBkRqkZ2SMU8UavUr6MrJ79cNd7QoLqslrWvL0jc5IU3R
xciBZgMUCxyVsYpqeA0V9zcs5ES6mAgZmr2p8uGYFt/NKmX5L5+/rxD6eGl0vp7aXBVsiCGo1IN5
Oe1XCNfwTBqdqy4IrvRpDmA3+Z3Z630suXwyDiSC3BW/JcAqGeirTLo3SmKtfo7QQtU6bsA91CrI
r+QelonEN448ls1FzbsJ2SXoDX3Ve8s212rQvGRAJpOxJjs5s8eJzJU4dP2/VgATOafCGgmX/Vi/
UlPrypoL7OzX7wXyZT60eNQsUmiBmaFEnNy7UOIN5L78wT/qcTzX/aZ/1SPcONhquNRIJQPOnULl
ARbqqJEeGwlqMaPNAwobT3j6Pj/E8yEPxDYCPo+CyTt5qTcN2oUlqZqxqUothMJL1e4OXcw069JP
3x1OeiZw11ZrYZ/7mhcXyfw+SUkzCw5QQxPCvk8E6c7dI6leph+lyDkcqo9t/4lfr4ZIqYZ8P90i
Av+D9ZEDpPZihh/Wui5tynQnB0M1j5v+Jv4q9KwSJNr2B54k5zzqKvATqRztWEazgBNsTxYTycj8
IymYpsyKuKn//WUCjyR0HnQJAIp+mbM9u1aQJO559ECpKlbL95q1A4G89AHNbOU6+O7S+iT34Nw5
BHKSTpqeOb7vZEYaZI5uuSPd767a7uSMUKKlPZnp0D1BsEHPqk02ejGo79UcIZ5R/UpyvGdAhMSB
wSWSXeVZVtzejsJd8klii6TzqgrEVvUchx6/VpG3qE0NqYHYMRhLafEcABROLtoW1iCpF51icglW
e51uXmALkhWjEGfBsvLT4fZA8OUHCUiMjYJZDbfd7CrXpxqpsLJu6S9wAPQfBlL89cEqo5yc5iMO
9/gdxTFg1LhSWiUF+G8AIMqn0FsF79Y4Zwuet1ybPXoyCAeEcz01iGci+6m3IJrUtz9Xlpc0JFog
HbW18Req8BbCZJKUqzugzuGvzuJEcK2pY3ne4ju1lyVi706mvLdp+zsKYNcMcQS+8cDsrWe5eXiD
W10JkQZ7tpmzHcwykslhAMl88bkWHUnzE1DcWty+ywXjgf2Qq5nfYkNmoMv/x7i/5QiubMWmebRw
s3/W/vxzdLkyYWMeMSCKqncbd86Bl/Us11dMOxdwzNAHZ49ndD8DXw83wgLpxIgwMpHdei23jJMP
R7zR8Kst8vloFPprqd0cghx3l1mff4xt5LVOIkH0UxYI1lLoBe83W1xXnV/mZBOK6/O5wBJLPsf/
XGpXvNtQTrYpDhG5zFpuu51int6k5y9K3Zi+DSMIqmGJpDV9QawY5I8hBSoyrZZ76WfHuWO3Gxoq
Kjg0zYATQJtud3XXbkXh22dHlV7gSZu2u2/iT1PkJjFi5yCxWaa9IIlg/JlfJ5og9Hq3VBmopTz/
ZUPHNkxpSY9Ak0mUed4kXJttJxDeZZQEIpFVpOKS6l6CGzktpNg6mN79sgnz/pX65ko7WG8CZMUI
WdCPHqjOq7vWn6lQavitXt/+pNOKI/E2HMTgPOkk/FJj5s1UgCHF3b7H6KFrxRA7C6aFhwK5z4Zt
XSWD5td0NIT0UEkhUPOA/GFvoncxql8flcR3vcicJ4kl50EuRUc+kxj7sgENYN+vQqEYczIE8R7Y
vcQdqsBXL8xgvHHwtbtHfmteEG47iLlJN+ELYpc7Ff3v8ecE6/2/trGYJl2KXVxOc+9W8NfiWpwP
HRpNOBd9RBBHOhKWIdNEcogD/UCRcNN/jgnvbxvvjrt4kQrKjdUAY5rw+pL53NxgFOxbxoNsV+/h
JmVH1IIO4qFlDa60yCjHYFn53kWrXG6XiqqO7btoLF3FPIcmGytyPBfO4aPOxb731KieDraM+kmR
mOGRX7fuOOAWv2CCexcNB0VgxNz2lWcqDdTcWVhXliOKZgfXX5j/Ew/bgHqI+IXfHeja/uUeIuWc
LdegBB5creuDs6K0n0FiVCxbRhgcP+J2/8MlLL7hHsk+EDOQOrbcpfCl3Dv34e4T1z2sqz9s17lp
ngULKcCGSmBEajO6uVzIP4cYqXOfcQC/Yy+G+5lyjoCXCQ3hjYI3l5W3LykwRvvy1mqX3SYfgxP0
mWW1Vjx+3w1axiufeCT9W6Z+DX4Q9AmAbQobdlEyBgXTPj0nl0V7yaMslCsqQ93Huu2coCYEbG5t
Mpzbfm1zaSTzqo9jwLMTL9XzS/UpZgOrfQbJWL5CJ/amS1EUveFnRRppI/0sjEFaVC0qVxJKe5BK
kYdvw65yzCjCpLUnPgc2egWhX+cvsS3IDxzNmVzDnQPYoDtwnf0wKhjrnqgyZ1wFnoxQKSUZvLhg
WCfWP2myrzJjzMHKzqmRAFKfsjo1TjnqFYQ/9z++HAJ1Av0E7hc5568FvAarKpuMOb2jELYXjTuu
9Jmsyb3tOi6IebRQ+8tNYMgXK83B/v/m+lNS3Pz4YegHNwHppdgbxfEqzw2U78NB3Z/XRYAx/Cj+
7ovYC3ZWNIn+Lp3OsjNxzPG9+jxktbz9Q7ar6nGyt3a3iei7tm/xFr/XPNS12UJJ2TxzSfsUY5jt
QwsCOIdmpimuv0ChQkEF7AuEFmGrMDBA3iLIC+vc9in3RxoZKCidxvQ2Gc440cSAgiAeAT31rebq
19pGFV1JPHx7CDOZEJyILwFEsCWs5MBo7oQRzUqXlDvjcFA0qxogqroN9WzWIBwiqQX5oV1UjVOG
y0jzD/f7ZklwokDVn0Osfq93/jm+XdDowJ8fM958bKryTAs51dIeLmUUJhqLTwBR9Rc5fhovVQKf
j2OpyhTpO8Wr9v+gbZKStfuv+kg6vzxJHWF6REmySfgeCGHuSwfy1+ruk/7Dtfqpplt7asF5d96J
X3XyG7stQsZpA/2gZcgp7rDntcs3fxXjN/dP6/UT8kh98X/vVMaXsEyNExQZrgApazDpzL5BNl40
T5AY7eEDvtwa74kgp5FTPLY20pmDZI6EMaqpb+fzZxNHYM10LxqnDdYd3wbXNvHN730qbD45vYGW
Zo2gRlfstCdqcE4VuN8kQkZjMDYaJ9/eSrTcPQrLw+EAliOav4ExxTk6w+LyhQZXcAeAo6tJGSKB
ZNfrecaO/IW0cuQ1TwfZFHZ1z1Vj4E/EataKthEV7YlBVUuaWvBKYyX2MQu8N8S1R4Q15vPJrhNo
uHQ36a1AbaSPKc8TZ0JrOB8+/tYABoHlc7U7Si8iustKcqDnOnPtrVqwlIcwFzpgweDqGs92jLkj
W4HGFMZDmQsbSQ7hQLJQiMvL9vSYAU+M4OJEN3b+M8yHrdz52htZfKqZPeTQplmdLi4W3Ko3wvwB
/erGwlB6J1D4XQhz/uYNQ4ch/LPHFjiaWt09Iixr2lYCAl9XQ5LKj/ap7oWQ5dKVgfOo77Zq0RyR
g25xq5QoLGJvC2isqs6BCezNNYr/lits5KZ/EbpoFs++/WchBtcbzOzvTUMj5PVi/Sv1cJXzAjWq
t5C1quLD3blSY41/nVNuaCbdkM33R0OIYat9xQ+RW6K4cEtHZqaVoQvNzsJ8W3cOpkDVqHkJuVRx
ivsCN67hqK9cHXaw1VV+rx6qBnW56opXUzYHh1SunEtjqsIy+XphOQltHAW2ZgmBFboPfw7zRocg
iUqrMaj2FhH96PyEAJqv6JNiATIFBb7VpCG33ThFos8sNtY/dhCg2bK2CJaMILHmJVbCPds31VOy
mbrZK7t0ehb5s+35npEf0e+mEADIDR6MAZ+DZNOnb5UK6hbf7wHksANDyM3quUDPiY6gCUFOePyl
OriLl9W+JxEgdTm/i1ShLJrKJ/8dgEGxjcCeL+M71p9S2godroYfFAGL7LW+pIluJPY5ubTJZ/hv
9EQ5H0DTAcE3X3f28fxI17mbP0XQ5B7grZKtU70la9iRxKqdEbeu51XlrrA9oK2NtmWKHIpE45K2
txhpy3rkjUsBp9CB9edsMgPJWIVdMEElHGL+eZpXSofkoB0esJE2sAEswzbbTBSCk6zUpBiJ3oga
1f1Y3XJYzIHLQ/OLAQV0ZNRlrTbZXCvHwppyYz0ERoWOZPTJNoA98IwLcXCzXEQw/x8OBTYDu9HZ
QmxHj8+8HKmBApAfUw2/NweRCwoW6wQSTN1AX+jPaHX3fFtvIgJrdmLePaPwoEDD30/j/5ra+whq
aSdsVlK8LKbdnb30CPw8h92jFJRlutQJVjyU3f57+bnrUbJXjmBjkxx5KyoQRIkPU+5C/v9N+CIp
Xd7GSMfX5xUGFAwm8tpircwtmIuagTyWy7ZQagbEls5pwgmracm7Kit1gi9hZtxuzlNEwa47HepP
lJ7C7HEnvPX8IuFZdPmbr+k3LZsmFhprRUJmmNvaPeDiYm6xeSav1chOuQT8sZk3iozSOhnQv4Ws
DC1/0fkWz5X8qFqSB7tZTWCtMwiv8JyPY5E9KjGrVRduNmVVmH+t4+YOzQw8k1ofYB9mqhZeLzxs
6uMgin7JpQRWJ1ZA+U/Y7Zvf/WAevzslikTPQyNLlfnEsw0wZC7AkjpLOXYSAbcR9YXY+xrNMb2u
Hv7mvrTy2pW41iL7GfKmEb21gsgQvzK5GzMc8tbxFJYGc1Ix2BZg9SP3HDiFMUZZJqPtdy/rtr7e
eqZG8bAKMVM7gQfbdhtobkDChmytsa35ma+aSKsLkKmegVMwcCo/bnQMfsvUIxPW/cy2RdhN1X/j
rznsHMq98bI62W04yV539p8aUmNXfXedH9HarRTFgmlAJpAeDtMd7M7Ih507Dtk/1iCdR4Asu0k1
AMHY/2x6lNqEOAtiqPIAWMe5j56Asp58QamhsymEl6Gzo+K5ZxKAa8OExUA/bEfGbwA2CFIymZf7
IouZCOijRpmGCL06Xe8HQ2IZ4XZYg4G/gvNJXzoTuHV2Ymh0wuCzlOQTtgUAjrLt6GUYouBIHmT7
uTcGAOvgdvV8yumq+c18ogfffbEo8SoN1eKzu13izeLNQu9UHT5jfxKMWxOkVUINM5fvh4ba3QPt
UsRUU2bFTsv9pkn0Q9ayy55uWZMUxRHstn+FBUypT3ZAw52lIbFb1ws9wJn1T03Am8sBpHe8gW5Y
GMizolk2Hak9b1yUR2QIy+YhOyl4AGtzjIyulDrOmQypRvu5cAkry3IR3suc169OREQ3RzvR+OXT
MKmd6ESZHy73XCrOMuFAAZ+exBnoW5ETTp4QEl+frGSotRUmb6iZbzdzzMiGkN9pp0A7M7fUgUMw
m7/4vG8yKbqPP+J3Fxtl7NvqWng5/KuLSKyesPNql7xRE9/vBK4UeHnJNKgo2BODDILuC1o1hleQ
mMI0/GDbViq7IhCzWq8QCzz5kFWAzFL5LVXIORl3hU4edMHKSxqN18KRDebzMGA5VlO3azuEhWko
kRmmait1c1E0MgoEKlXaN0o7azg8WWxywQ8mOAuOwv66fPeb6ZibkK3wQywnLG/AncVW5wHPyJH5
HdizlplWBY/3QB8z8z+/UPMJ5t5UxeUyFN2TlVN8g1LOiGRqrzlbguGwTk7EHzeMIYTbLYFwz+Iw
xnjJRF737yS5qK2dXCwgxt6cA11ewOMTlDLxoXvopB0fWKJVrxK+zxZRkoron+KhPEWStN8w9iGk
2Han1pi8z8wE9FHL0vopwM9oQrxtHrq7+jORpT2vLhoG5XcOnzeckdjJyd6XoakMo+W04sM+QsTb
kPElegcgZMkvh8Hp5aLkdQScUAaQM8GrhC07vWgz9so4nDRxfcT3nwozAFmt8sCRM3atix2pMsdz
SZ2vAmDmdmFwnJhi8TQYI900SNiItkwjS7Ru9fE7agWcP9hyL0GKRIsrV/2Z/FxphJskP4cqpWhd
Y50Q5jbbeHr4YwSLokuHM20wj7pN3e1IHRw31Dy4uxieBXWzIRl3DE7FR/hXbZHNWjHgBGUAEwV6
dBFFhgMRxm9lgrSttlxTjFYJ29hNV+mfiHdQKAQVMcZ9VTDj+PbSFiALGW9qCazCPoucSIsw8Iie
izAdOFKHT4b5JNvfg1k66yxyFGJDtIKxTg2W5kdmZyl6YdiP1YpAXn9lslYmMb8VSRDnzuO5qEym
GKxVobj1yHfHVNSGnP8yXb/Rpssjaui3Q3A0J9Swl9kLLP/8F4GFfPGBRC0nt/nUdS7P+i65Gpft
UIpEywfWTFp6ZbPWUohjXSuRJnLeXVD1oDKHmrkbqZPcPFpTX5MTpTuw5FKReE4zu5ygfFgeJazf
br+X1hVIbXmmNx1+NxBoVRyhGjf/JIFC51hiKilU6zqU8eaZuZk5z1LxS9M+KmP485HOzZFV4q+P
8Op4Ww4h4g8i7B+3diw9rDVEq4WPbQDLNDzBC+JE9A4J9PWpnmcE7IZy7b72XK4zzMi3uv8xhQiq
ntKrA/ZFs8a36LAsd4YnYW70P+Yq8DXkXwCCQEP3q6tHxZd2j68EyJ1P0O1azPYy4m00QMFJ1B56
bk/uGYDYsJHfIp2BLn7LMJrOBP5t0A8/xRaMy5woj317f/C221gWdW0QgGVD+Dpley0zUJhoF/Zo
TY09EZTvf9DTq/TGg3n2e2cvF8K4Xj7525GBmlkyKS5zz685Iu8A9uljVPRcDPPKJ0bKTIYBCV2e
ay99xRSiEB31UhLSBP6E3FKM7Yz05zLTeUw9WxgmUdrZm9baes8MkzOFSyB/VJKcSmFIOcEgei7Q
q2hBPb8QKNqw6DSVB2zKjulIrV3ZrgdOkULf6rBVezkrBl1jmStRIo2jl+0xVSuZoSVH8Ev//ukU
24EgZQW7YM1Yv8g6MmDjvODfACcrxrzm+rvzLaFqKtwCxejqGkd/GzLYpIm/OVK33Oio6ub6nbD0
20t2xGayP9ycX0cjMCFyQj8mRjSD+cb20XPkH/ltDMrZAW9M5BTBkbFrcbLZ+PvYnSUMpn3SB+/K
IEhUKIpd9ev7ZEHxai4ZUMSJfNu5dAOJnqJoSyk5/c1Z2pMca1npmezhrFZLwwMVh4XdelFHVi9h
UPjmUXWh9pBSowei9TfXLnR9si/rfbm0aX2pTs0GWA02CmWVB4cT9DXe4cLU+Iy/9F63jcMwUavu
t1+1HrAMNCQKU+nXbHZOt1lddULBpvXTZ0OEW487dw+TOxYTBHyDMzbKsYlz+3LqSUejMip+NzXX
QKtDjqtyOD2IZsChb7WsiJ1KbRXzbcznuOL0RZ/QgkeCzO/zwLYzlhfmQg5w/lX793s65m9x55kX
7gUFDaP3woJGPnZ+4muopXmZsMWBGUFSdC1BnVKXr+V8kqGWRVwAj4MzR54u4sykycLR9lATVjN9
bFV5+ROFi9OvLes3b5YqsDJn4l9zgfadmvQx/ZH1hhDLoQ1k0TrgJ2b4kz28R+lya2NIcXnNOaLu
54SJbnyXw76tms6Zo9dOqrarpi+cIdEw/vBhViG6TPiZxHyLGYG3tp22gwA2o67ZB2NgERoZTt4H
7Ykdsq597TAc1EC4jBW3CVygAa+xRW5ywZ40/mVsXyGROCcpLGev1z+HL/gFdoNpT630Up08e20g
tzFPkW/hUWDxocMY6DwKoAT91YAo9Oz/fm4M9eagk65tljLzjq9Kkzfj6/XtnPe8EMahw4JOloJG
BUSgX+JuBoeloJX+ceF1Mod2Y8VlCo8CtqzNa8tLwOvQUMECa49e/P04YCY01wIlTvlJmhl5p6mF
XebpbH3W5DGyioyHnj51SwV6t7HxxuOzXXCt7q5TsW+qxuTIamcnN+kA7wFBl6HXwK6h543qAzzi
TLb3aFoGZIzIQXZ33Duu3hPMPvTKqXQg0x1jKGf9FKU4tNeSyxADbdt60kjlX30+bhd/rodaWNlS
kegwklk1tW0ThlEz4y7iR/tWfKCAbIbAisSpSdUdXY2Nr0Z9n7+vWF4sB83RNdlf9bSZett4FvwY
vzUPIBNfH2orZk8LJnWVgOpOOxZkXYmOb8cpTDHi8EwwkQzLrRLoFB0XXNpmYdQwxGHWVe81se7M
8ERmOlO6p+nezZRfXJ4N34iTNjkuh5lz3p3sPz2GCBGEW3il0k0T3mnktCgOLkrLcm9o/VlhnWAA
83kaqJIEuK+O4nL8VpJLYnlEYrhEfQTQXgU0TaMDv6G/viLl1lmGMhy1xkuPTCHyEIS5qbdLy+D2
Gs99lz6eCtZQYWph9NrtzlSgqzycRX1npFgQ5ql02+hX067krHYRiBu4OvWDki6RP/MR+Doz8Wbi
1qP5iLcAqXS495tARtfijfT7KnqRFaTxnB6eR5vPIRJujqGdhne6Rq5soTGiVRe6XcScq4lWzwze
P8sc0YbJdkgWzPwpNIyiMcpg9ilqfMqoUqlg9PtNjZsofisQr9wYYuMWFBsZIIxjEYzlc+ExeLOV
wo1kbFcxosniB5++Rqn3tVR5+w9XskKoe2jEdgYUpiZBPCsMkb6ZAaWE0QCKsLXRmimLDbaVqw09
t7+sgh5XhgyKulqdbA7578zld9AWkiPAN24UiNraF0OBsgU3x3hQQ1fjFjqA+CnuHvkknWcbeLxf
BVpd+x+WVI5clb+HsAI9tAFZY9tWhVzvsba1/AKEbczeHxCAFZDXisFssafXm3OrIjfY2wFbVCCB
rSLNLw3Oi5iMEd0RIatM127IiOp4dZ2Sg+A4XcVDqo8milonF5kXPHh+rLoONTOff+Pk+mg04TXb
z+87WUrmFnBFoi5TxOMMjDzqW/drI9FeGuI/ha62ZEQfngvHAt+z7+ZROhagtUAPshW8ncxYUZKF
ycx69uuZ+2bAPG6c7VkugU/IMgqwU4kJtSaIuUgXYLwCS4KrG+WHvwlg6GTHE19jn3Nv+x9/bWMe
k2Vfs7hwGTEnmYvYCUjjBkMCWHN6QFaGWMlOCBIaequMaXZz8aBKEd8hoaWp46S6WmQnX0NqN7WV
Vil/VgRMZKvSjUshUHQ3TFmpHY4iXbRErsJ/p/DCYv/dz0rMCPYdnVQvSf+Hu1u3DCNm/YelT/uE
HmPnCDRquPsxZ4Ahg0W9NVdYjEbuEt5PeZVJ2tt0Ic/jjJ1ifpNNhOAKNIpFOooJOkO9YZ53/1Jf
roXloyChE7IxRsk5rWfuq6a0P7UlkgMDRefXC0hsFHhjW+TOSNDZrfqgoRBbSs/nRiijqTh19w1R
WAPMzthmKVgjQ0AfKkNsAm6Ovili5NAtffpfYemlXP6UdOTUCqcP81zRo56UU2wmc+WfmuoIOrOT
eHgRDHiJcU5Fvot5iMFukB69Dp+EhAHiV19vQlR0WP1wI3s7Ujezal0kzWDQESFzzIh2YSPE60T7
5Ypcpv5bBdEoXLuLK9wncxrGhMEL2kelV58NlJ22jfOgHNxLcnnwM6epdbTZwN8aE63XcTVOdD88
a6GFUSloxe5uHRLBqhU1LDn+TN0B/SmWXbO8LaFMo3MzTttXTsckZvJzHNAUpZ1ughr99YggK3a/
gqJL+3RedZGzTaCefczVSzS246xinhKoytC8usejyZ8X1T5JAiQ/h9LNyxG7ZiMnC/QggkGrib5x
FnTTUHEZxQwKMaLQhWDHZE09F/ieyS+qTbkLGJaOZEdFeR21jwtOBEOo1fnSnVEZqZJkZY/FKZZ7
059t6UQNcFsse12SqmJMxhvTI0rpO4wMnfyDk/C4dycN5aeKEVc56PPTsDmOUvIOD2bvuxdaOA4u
o0oTzJgwU8Ak7XZDuxJA188WaoxlTT3CB+vWxcT8nyJ4BCuYGOrVwdn8BzI39jcORO6l5mmdu7v/
8iskpCKVwQAj32Ao5eFyF3vlOBZhKmjU3d2UQeNQIwGJ8d9J01zWMTHfORJ0hxCOpRYikSGDTzDn
g3cKoNjA81GGmBqqLpimYftAfPrhRBsY+j5cz7p/4ymgLgvQNti0EGZuiiw9oHGDCDBRRh89T3x/
ZaOIBMRA9pguvhyDKulQBsaxxTbnPq5jU6feTcaPRYYNxYETEPY5Hmzbsv86iwpdVKjCxjwy/7s+
FGMbeMMKosrILqoCthK2EkupdjjvpucyJIzXcD2IgdSJKVdZcEhy81Dxj0gnXLQl5d9Dcw3zhXYX
FU1NoGiRBL4OW/flG9WxZ1yujkoVhMaSSlL7zY2KjnhJFqvJRbXbhrKEFI+HSVGolqKhM53iw6ES
j47obnu4MrD9p/E1O8T4H6EJZJBzJnEyEYc7ji+mf4kjS/sYSSM8V4eaayaEP0DrBVfRYpXXQp8b
Zeg2hRzu9uh1g4Jup+BjtIChqwkuugtlWR/E2Vt2ywsBM+mfyuHBU4nMPe2ZcryY8PGge0hKHBKo
6qAQIYp6WKD3Lm3MsZjBF+iOyxFIAWawZaBCSCFGxk7xpGzKYH39qls/C7nAQRQlcXlGFq3+glCp
FoWYnd8IBLQeAkTcXdsWxYKWRrmytrpYjUcS8pMFjQDdQkv/ULh8VT5EmcmPLEdcKnIKBSHmuRr4
+RKqLD+tTFOfhXUPSj/NS1hBhxNJmgHsccftVSC5u6EAhgC5aVx5FHg4h8YiCInGUdqFnrITA/d+
2q0Ma+HwbAkbnwetbq4zsw6uTsHyvUwsE0GbzGSaoSfVl5tZIMv+SwjhGBp00tGukPWfy+Ig+2yI
7EksenzM6XGTYVilkqAi8DXFJcMKoY3RnV9DjS0gneal3VjMepxHTIdicOPbzjaqhe3Sfx/9XIZa
ke8Fw52AvbAn/UpTH23NgDJDXhESHqPkkEQxkaUDcWTBSrmcPyQ2Ky8iO3x32d6vYVQGYTdOJopT
MhDuOEr/OUjBRmLqxN1sR4RekWu6NLnXCJXlfJh/Tx/YshZzYA85Ertp6tjqzeayQXZpw0LKoqgn
x5Bki3ghf0XKG5t89S1MPQl1XujcebhfNoDMFH7eav54u1r1SFBq25sxmr4DRkl3uPVz7Og/soBN
jZbeCqj8ME8ucPwnfc7ECPZTeG6WKRku/SltJZyokYBq1T0djcphrbAdRF52ldNTOoT9Vu0sNZkC
WvfpBJ4Cs9k7bOGn/cTNDNEpNbLotN138arJ130owX7UqE+cdqgm+HP4fuFa0Da3fxQVrYqvnwpP
sOnHArrEfIP9BGP97kfQWowjzWVNAKt6ggSV9pB5HyJqNxSgNphPksH8zB1pEyEBq7dFzSgivI3+
InvQAaHCTioW8O1Ig2qRT72NHNga9VgOPwuWL5MadX63ewJRucfy7P1+x+cOuCdjw3RzLn+3NkST
KobRVrX8swAS2lT/2VA1/YTe01yUzClMtAxmiRCzHhIMGFNtrqONXWsXdOdGvn8zbfb0mDEEMc/u
+jXT2lgpEUkSYtQYqtoaXd7vPc9INntsgvmqiXZ5KxnVS5P5Skl9stL73qWWPpLcxELGou53549r
rZUbDtG28uOhoonstWYtkTZq2HFXYBKi9cUmL+bOqgiKWrA1yYnbNviP0mwJ1I02pd/HN/SpQ5qw
IJpR9wUdIkbbMsV7s1riXq5iCRHv4RN3gEqPTq+NABXKGT67giQM5Fp5Nx/Bv+l6sqDKXX2U2ma9
irtxuoahNRiWm6l5ixVN6PV14F4QjCtLH0yQRpUHDzRc1lz22TYNQ5//k8Sm/+Xfg7oNceG7n8pD
w3EA9yUQmYtcnHMEPalm7cRFgkOsdn7plhQYnJILkt2PwkY0SAAqytccRWqOsLaAwvYedtLYm1JS
+xmdG7KJW4pMtkl10BhVAsBwRbPiXNwMeEaf8fpSbFpHxKjWupqerwzc7gmYRBpBT1/hXiFl/Uew
qgxXPsqp6ILWSX1IQ+0GbuN6miav5bUYn3slpiMGQLUMRpIjjE26QdwMzLiLAxIgq9E1N3zXQKV1
fp/ITzFxoSxWWNkoZHPiq/5NqmdQQUq+qlU8dAd4vomFEy4zMnJs7esfObUMAvOX5zKbwpv2kRMW
TGSAo+Z/TyHvTTDzifBqjJtpJv3KywBW2UXz7buYi+EtOt/HXY5Ub/NBuc0aX81CYF3U3BzcePTz
2LbOm1zcuSrY8SuEpRd0NmbIL9/6s78Uphb+vn6+0LLjfEtDwQw3Ny8D5kGJiRiR/o93ImkloQbF
lK+tGV4a6oEov3Ih6K/+q+VXxXlllDZHrqSdCR9C8R1xKWG7CtwnXmKYDxFtkdD04Ncz4n2GrfTu
QHX5S0BgfPiCB3nCAo6lKnqC2mh21L5hCY/+jvStCaPdahVbfSevGo1mkTuFAUi6UY1oONJNE6oW
ViqQ62UugDRHXsUURyX/3U/HIpfufF2a93eQMasnBzqCd0r/mx9BNmQzPRCbUSEmJapcgIumtqqB
Ej/RcjXDQQO31As/MEtANbuDhEHehdJHHbud6hw6ayqW7aOk8DPH+InKkkSKVSXD5E2cTg/33TwX
IFD2l2Ig9rjy9O44ED1qTxWgNDLrD8lwFQk2vaXSuJ961OImD7ONqTknWp3Kze9XPPBsZG9YNBJL
WkgABg6drN5qpNUrwF1E7UgPZkGWINzmEx/eawHScXP85Y2V0j686M8rh/rUD7OKKcozCAb4AKK/
KkJpILK/vh3F7Gm8LAIdXXi0LTlDMChQJjMxFGNThNtPS2LM2RtAXoEkWGI6ZfWpmC26DDJJFzxg
BHP3zRskv5l1KVRDkkxb4swxdZXRU7lfWvHqvnmTvw188HC10QICvKnGljRYfXEFnm8dLX0w3ySG
AW8l+xguF3Ff9QTCxyAAHWSHav3o5nVcSyzrDcd9oee4PRaEOs5hx59XoYOFPjJbCH2Yl6dfAJPw
3OUCYvhMFqYtbbvi66kr7lmUnLG5u/kS67bdjPVh/G7eEUkYyysxCTx080Jf2E4n2fYX/YbNl3Rc
/luou82hfDf9KwqPpyhdetACMh2fVWUIloJa/cT5uyHzi05lAMZlxr3ZIE2TBJ4eAn+Y7m7ipaRp
r2qvdKjxFFfrm3IETxT4AAheLLbIqQoHyQdrO+x62jQsyqD/EazydtkNwgwnK9dW+YkZlxaltgNH
RbpSsjvgd4Utm3ZnU/zIEpyKNqUPUJ+84cwyqSKFadeoKhxM0q7Wwe51vyhSi/k7tlACdNu7t6fl
OpWBye3cV8+NxPlv50om6odk7TboX9z/XtDnu8fUya8SWr/BJZlKAqilKwFmAEpK3OkDC7qRtPOC
efdzrgtou/qpMPY719blj79Me7h9L6jDrElu+uVG+loh7Pog0lGbhLGoAX+ihmmn3BKtS6t3aFDb
jRW93zZJM+rDluBYLJ2QTEqGnbKlMoFzRplESq333+f3GXrOhdUnrT+/vjNReZf/5fn01Qwl/0Af
XKj+bycL/dAVQMHsOJ4pGsnGM0amMD/D/I6aZTMJ3lp47RgqsXwUaALHhuuFMOsgQiNVEFjT4qbM
U/4nkBODOXxl3mPqAqTRGFd61DODrtTVlhgCkK1OYGQrZbmvk087/313fyEdDFKzWkz8nDcZGBX7
U6btJ+ci1ognrLVcnw5tJyyFciuYW4CUal6FEqcTgIkwLNLABpVEyRGNQGOi+SLpG1bK2kAVa3oV
oh8ErP9OoTNd1qRtorqYCm+kQS/Z1ClgXPgDoi4IaM+296eCg4k2+4ziYf62dmt7fseeX99eUL1t
yx6SbNYeDoOxKKKVSMjXfqcedzDRNphojWNvZ3fhJIEnTnA0mSCZK8eHb5bnBQEg2LVlW3qBeEOH
NlEu/VCsA9Sw/ked9cxNjJWjG0HftGqL4lzuoJk598DSuNCl6/JZesyck/bc5j8marBkiLQr53oU
guwSW5DKNO56vFXO4PBGqqNdiSTREynGJOZRLTY6NKtiYJr9cJrcDcJYxINwz5AysT4ytefjg4ip
Cavesv7rQqamiCuLlod3kyMdFQ3XCPn6ovKBGnzU67UgDOfkSSYvGrUoPuUNU+wi8lFj0wAkX3bk
tsfa1FiibhImeMzunbtc5eDmvtQTcGN/ZYfCDvnRLs++33pbRFaO58rWvE6pk7cN+rrK0gTXdrZR
4fPtogIaXBmbWwCsS6U2fq20xHZm6p/EgcnTOWN6j9OX4T7Q+ncRCjCoYkdM7BlKlktsACWL66cK
o4SNYsgSvi0fcV+KRjjItczzvybFkIGxQQCVAff/oW91NCzqBbVpieNvVwlRUnv+s/62inQqEDrQ
fzjH8iQVhK7jTU+jUJArZaZhN9vexj+ouMtPQl1hwo8/Z+skyiCYXgMYv+InOIzcpqqPI0UPyZsG
O/WfZZWeDL7YC+AkQ4owF+AJzqH+r5lrfbTgyEjMBL7PDrK9Pb6Z8EjpLcvnMu2X3N7DChz9Du9T
EkG/BcK3xSOfzo5Boy7ma8GUJQ0VPyxonVuY3/fF/TyZTTdSM1ZsqlFmYYpilisDj34bwY2uePAr
OMNKa7Hdtaj7Lipxdy/eFAdCFnDMJa2iSJEUZ6iFPmkHk3P/wc5q8Mzuo9EKIODBQhavTLxU5zml
X3wn90UrPaz3rWIqWMYs16nl6JJCkkLhR+6lsfqp2VHMDAKL1JFdFujaUU6HbcZLlZw+sC9IrN80
AJZL7iX/yqQjNvb8zeQdyA+h1F8LaCIOuZIH4MpyQCyIBBbzeDbf9j/5S6I+JO0i96cJBhkJsw74
bFQ9X9fTvCpEZ19OjY4ZCX0ZYvYq43oboF8z4g7vxFyxSLz0g4EAwbWvvgCcZtB8qlyxEFPpZPIi
2Vn70oCT/XU880Hz8eW2GdMZoEI5kTJMO6haLr0b9AK5q/AKBhxzXRcZSNbHmOedR0ApQt76tpsW
mEI2gb6ylGSe2XTRXI7kY0R535qKHlP9Jwzrt8WUbjWUyw2g/H+p9ozChFXCRAXA2NzHCzKdFM8Q
EAE24ItGo15bax++ezVuP/NK/w9nwpf4rlgdAq+g4FmpRCQFntHox0a1caRQJFUrkR7zXDRGSytg
Z4k35RENTbbtxa62v/TT2nBx7O12QpeG+Bj0HmFlToVCPXRyExkliS/QnuA27KQuQGeDglo3gzqQ
/hgFjXh6jfZMWRcX1zR3MlSMJ6qDnt/EWlLwZE8mBrn/XImV0Nnpdp5htzsP+DOFnBOamq2Ks4v6
JnOv4N/JzhX4k4Wgqz5bTZJ6JlZMZfv/bUJ651N4NCIGdRPM4LarXPoNcbWwmDWd5bBdwjjCIwk/
BGoD6lU5Y222vY/F3HMcFn0nLGI7XfpjEeYOEy8ONxexaf1SvxckIYMnJ9QSHr05PuLydGlnYb5o
lmnC09v6rRX9fgcrVsIwn8hORfnaLFyNYHX1i+BJtPcuc6Ym0UW9Mfk6kYwsdikQd0D3gcKTTeUk
yIfI1LOWcNXqGOOxfKmuhfkKOEAaPK9NWq1o1z88Wlbv0WyxT493pDjS+WKWKOQvmnnBvn7h9CAg
EDtFvj64vOF5P8J4PIWzPv628DOZLTuMw+wtAz5c9/3fHYR+xXXB0DaDgkPvfyn9hpEg+vLsOPH7
n0kQgovuiJY3MFpHVQxLvNiZ27zW5RPGrL+iADz8C3TIi/9veil8ePTX8lZH7v4ocdd1nyHbAiX0
x9L6NgMiedZhfbofZKpXThdxCl5m08SopgUGfu8jIex670ld59tvG++wGlpKcEcwlXutc49VYGjP
jKKJnB47OZ7c73hmUnw1jaT5KxX+Q9FyjjxMx8oKV6aXbtZ/8OBfs98OcoWRnRDMjnum+u2Mfizn
sVjyJrxNJrNgkjUeSjiuWk5lwK9CNIN5sEeCSwgaW6hJ0aKC441Vh6tkaoBEXE3IG3s30QXWZuBm
yVNGJfQqxACFtJheyud7GZ4hpZSB7eiMjw+tfiDYs/40R2nbGuGMtwLD0qD3AwACBHwTSy9cSr7z
cvgif7vMiQgn7mObMM48BSV2UxeU7pRlN08NNTXcgpm8J++B/4JyyngE7009GA64Jyn7CD6GDkGE
iXOucyNrRI4Iq8NbAOexu36oDO7/zTSly+MqLQdLEAFfmL8/XSVtG5BpFDoZ+ka95AIoMpJ5iE0w
xWOT/tfm0i5AEb3hZyrh/gCkf90d9rOiWl36Mq4wf2PR2WvdqxMt0UPsoCy+1F1ujj1oGv3IvbNn
QaqcyYxNpHaUXh5K4WEHbO31AjUqm1+cuEugb/R4lALDAGtcghqdhjq1m9qXJuTIPeQDCPsTntVW
/5omg0jTLN6TjGaUSxmtf6aIzLRR4jgfo6GoUTQsIYGgcDd+Q4P1gYllp/Fs4RFK+R0s5jhoB15s
A+BYZoP6TVCAkTdA+MZNkJAUpXLf51Pu20Ac20VOVh1B3DMRq3P20j5P+h5WmEHPVZo+9EbGZ1No
J0j8AqOgLZsy4eMTrnbCEaG9HkERvyX5EgK0gpswUEIBh6Y9CWZrc2dYwE9cnDkP3DKPUDIwynDb
LksZSMdgmPfpLQf4b7Xgw83zGlSfV2ou+i+UUBajWKVOt0KfCkeibxAR4+OkXltg5fVWX9K/MgZl
RQiqnwtWsdhW5KCYNH7vVdzi3aLRCD7EU6C8cmqLuZwDoKDVcWVqAYQ5kIxvgbMGhX+SEIWX3IZA
VApRq11SsSm4JbIPKXyaXJsLPqpaI9w8GdYpukVKIa+0r2MPj7P2j8FrpfxpTO1yFjUJu4vKR5V5
4rtYsbXqiHiDcOk7jT1sNvaRq5uKPAc7joaybV61oPum11t4xFjKmr0EC1CTLS+drfaWrNlMkLum
Zdu4EjwoREyS8PeLEa9tiSqYa4JYOXzCC0v4KAf4cfIRdwUDQ55G1/F5Y5cqZ6Qa1E1WOTlS5Jra
UnGbjHPs5scljAaHrclWxcOlMtcWiiD2e3BiGGiRAroBNm8BHh+EomdH4uB3ZK42TQFSYMWUQqc6
NbsHnXs8pPZ62dlkKxd7Vjb51y+OBVZHq83uf4aDknGhWZeW1hmV9iL0G3XyvN9jc9Zc2g6T2eQh
gark6XO3VoaRuw4FJtazRiE0o7WhUyRGKOUwsOwQerdS2v9NCCyNOGlrhdwJNIM32e8HIMBDdbtZ
IB8jCn1zIw38W9TzJQh5FH8n/w4TEwW9lysjnn9AAvCqAyt0v9o+0LX1UcMg1cuoIsALw4EGMU+z
GoWvGIXidQjdx3GVN+H3t4GgO4R1/D4GP2fECPwVyKpWOhEEwqIn8u6GZxmKSeDR8jqxehYHQLUH
MpY1lUiLNG16UbgefW0YOkrG6YOcgUF5h0KmmdzdVlRxS77boiBrUwHlRjkLIEupKup5p8400Hsa
uTXVvUM0gN26uOwBg5sAZBSBgIKYOkt3mWRzNBzZj8cF/6rpCvNvvGO8E7xzfAjMexPTZcga1XRA
yylyVpXevcqPpPlgctL2gpU/X24fmoQpP8dwxBsoPTnLEN/pnpRCATsFlSnN9v1WVDc/vvsQRZmV
Enmanv/zh+Rv1XXu681vURX6x2YrZ2VoYuZLa7hZCmJgvN/ip2OsisK24Z24ryXPw8ElKBXAjti8
uLiHSPkYNTSM5EdR9UioaNmRR7Q7N+Ps4s8WCNHtLn4HEe/+6mXk5v+g2N8yu2AHi3AuFK+xX3Lg
fHrnPANe4EX8wgC37dw3auM2NFDboW5AfhdT2NjGfgvNol8uvA9MqSquU/7FGmNxx6pddG5JLXQa
h+rB1vzsmViK2zJzRmqh0M/YYu4agJSvKRv1wMH2Y+iSOyDbcC3li0N19lqruPkrcS0y5QG3R6DQ
0gSoDx/2+TEtvUskiYv/PYJRkb5Nn0dX4kUDIrTSZnKehhfkHoLa61ECylKnmH5MdWc54TzF1wJR
8AosWf9+c4n/jm4r1zdf4fDmdHMwDlDmPkEx+xgcvZlLdWZr1ez2wo2ATucjfpLanQ5Dk4bk9G1u
hqm6RCyg6KcpsWhDvjBCgj342py88Nryqjwx7cZGPnLmsZqlw1j9ODwSY8dmhAX49v4p0Tubsu49
8ruYJXDnzvEDute4rEkfzV/c+kT4zBKzzhKkbSXGPJS+7RsJa7+1r9twCmc324RUD4tcQCtFsJEk
au++X+Ca9X/FDxfGY5/riEyg51Yj6mV0pDbDqxckigf+o3v8ZHRRpT10ip7A16ZIsND2XHk+qW1f
J+syeagu6PknfM2FEmdxB9RcUtGn90WfbeO+otdixPNWrAzLFKACtfamxJdPblD6Qrx7aHtXYHie
EKJz7pLBleKJjOPyQ52cw1lAbpIzyXT4c564DlVc/IICb7s1kk5Q36xHVkzD90A1VqfSijxo04/H
E8aMIKamhEHg+QmA3gh/pj68XLlp6XXuosMSM3r3WSgq5BhFq6o9rfNcERPocIWwvmqPV0YkowPy
ASA992ljb5wmD88FpJzmlUvdRAbLGYMkeoDvZl2E48vPXTHfiUkr0ULZQ4WCTJ4jJK4ry3zibnbh
qlytxoT0syq74WnS6ZxEnDXxVyUfy2Aw3tYOnyoa4HBoo3tCvqNu5MIkFhcq7IcITfuV48L6+VcZ
N/OvVJkcNiO55chfcUKjPp3DF2006sEISWq02UDvQY7SbAa5qc3pmGuq0ou6cjxYUw10M2RTS6ks
hC6IpY6DFBEygHFQwJqLfi5v9x6hTlXwN8NaI2vSlaUIS/39X3lRO2I+OzBiLbhLi2mF/2MWWuCL
JE5W2y1pBVTKW8/MF4WFZtlZK76qkJ7Zkx+mHUjaH8kNu7olmXMIi5gaQV/V96BvxbutxXGuqOph
nVrLSX8tYyPqBUzP2vBCM/PpV6AdursVxWsOAyVeJI8mT9cEk+EU6FtfXf6F1nUcXYoV1GN6pI33
ScVYHIlQpZehemMCg6XsnFHj9AevSRR+f4mMCqlH60r6gq/oShY1PB+uwBCrwqwPgHdFb9yumYe6
WlbD05UMCYspUgi3sooofAPkzfiyFiptMT3MVxUq7PLtjselHEUz4DOmyhR3IrtwGbIfh398lWyC
wA6VDrmZ5KGa+4x0ktInO59XgTp9aS2DxhN9aq1hGUXQASIYROB16jt0gElfGXOo+7GOanYjAARV
FWshUBUpb4RgtJPOg2kab+tXzpJtaXZxJNxAIM+EJEUWznXft+eRpAra7MHjuhcwzyGnM0d5ZasP
CLYUQUmHCroHhCy4texUF5Oy75O2HbG+wXv4XfXkNTsWGsqGbrgBTQBl98UK4t9FvtRp4D3CfH1o
UBCN7zXiFlSGSRrR2ObPlyVpwv2uvWI3i9ykuMFnwUbgXqrm3Usob7Zd7UXv71LDau6Ppb+qEFHP
MM2m9KE9T8eH4ejRqoRtGENUZtIBV5GlI27DOn3jbiyQN47Vqtt3mzRJIFKDSGosRDo9Xh1df+eh
D8aSIFvzv+MswfBF4yNCqVkng5M+dRI2I9b61xj8CFqK6QJtGCM21qvg80qhhqk+jntpLNOg8/JQ
anaHR4QBZxHiMdlJgY9VMks1cMVAeO4KYfPkJAPgriOk3TKRkSr43GkTsAgqrDamgfbkqKbPHmcW
aEX5MoiRI/l0BB4UQzTC/5TymT0PJWCNn6/oIcWaZ/s9n0P4vp4lVnDAD/iOvCJPWKsCc04/pPzm
ZmYma1yq6doVyur2qpYKyLkw2EbNBh4rMn75QPrnWJQQ2vUtQTU+3gXriWGMEQ9Il+27lpE4rdiA
yPW48FsI7t2+wQsSa8G7VOsKesApFmcKj0OBxm6o825aqW2gG2pFa8D8V5BdeT/Jw6h1IVl0HDiO
ekYqx5EQ0eK9ZWgfWDUJeqSJk8PrnNemWiXYLoQQCDgXx55IW/cA4a0z7fPjlfGOqBtov0VJXLqx
v57Wu1Hgak+6VEAyujPgFK5lntfTAwj0o9P/R7FZJcIR8b5152bLT2N92NXVrdfYp4SaCaILgJTy
FP9LoQzTPLaR93U8VfVh1QsMiT+72cuVLaFJEzj6D3IeovFGYwkZoeRJILbfQ5jw2JXPPNpzPqwY
QnQ0j1ybU+M0xiDKKZhFZQG7GoyEnJNSD5TUDGO9EpkyEfGJ4UH0TzWq2S8E1GVWQsKXnQlSNntJ
NK379HmHP9/SMCO3FXZqxTeg3FDFg1vdyTrEZtquf16XiZp0ob4tk2CGDIsw+Flgqo1ZjD57po9P
rZW8F6aJ56Fwt9SRcB2pXda5Rz7uIMP/MEmZsH93J5zo2hW9yQ2HQCplFb5IpuZjQkZml3y3zobB
U6VNFAJC3PzH+QpHf1sHJLLHjn/2LNaPWYClJl49uDDGI0N41HAFOp4R2yogj1+rKzTpNvXH3OlT
pGHeqdmVKdxJB3lH6NzivDRZrocr2d7QprKeLInqpN+ptAInAWkIYUcSxTE5kLpahuF9CqVmXM0E
39qt/66p/oOXPCzR9Z93N69nmsVk/0ptmzHwmWiBH6TsNfKqzOscOTKj5z7aNliImcyprZmr1jFr
qXg1NUgMVF6bV7H8KMe2dsN+kHpGa1PkEGq49QkSxZ8aTkeCjXUkbgKSP3F6inKe7II938MyfCie
7HJAKThZREK//y0aqT5BuORL546p9bJMVAz5Hzt1VjF25b/2gVoln/6TFdT/pybZvwRbI+fYWIg3
7D/9HXtQEbXfMd/QEytapg69tSABeT0i+bnKPxv0sCKhuVeXjv7UsSHtScqi8+rw10nWgq78nux0
ApZPE1bWOVwg3aSHF5IhRXPPOG0lCQaUSTTyXDZVq+ZPRp5AU5QCtl1zT2XdS2/RyULLXB0C49Ap
tq0RCooay4V5kLTnoMFgH+uaDiJ4YRVK9J5EsS9Wt+gEtE7g3oR1UnebF/VnEPxN34Pn4YejLBMC
xqafs9IvS37DQ58+CYmIyO05/QqJCljxgDP4QTn3CNlNb5dF8280WR1oHcXLDkEtbffYOoGmfIJY
+M4WZmyxgCeGOWJ15s42GN9dYiSQrJLUZHc77jlM3t/QzzXRUs8b6A/HexnJsxQy9QgHhBiOYIvY
8JL1eB/tXYivYyhCvbpS4oINS8Z23QZgX+TcKRf7W/y1ZApwZtXwVJcZPT2bBmX6fZzPoLe0Ois9
rsVqkAwozWonGW8HhwvrMV1Rf/9MsI7Rr9kKXK/EdUzxuED8mi9rDXq8CJyofMg6hywl8A2CQwV2
DDX6CHUVKhuP/mQ3+TAjLDdUdX5HKjinkUo/T5zqxz66YN/A3yOY6Y8MjPdAe2w90KVzKmypSV5y
xBLMjWlJiU15+8DawKOcuL8Oj8eU4ZM0S/VzbLwr7v6T+xzRXOWSQrqy8tUN5fw9bkUFCp5L6Enf
vCpRS5N+LWKW1CXK4kmDhZWCxkWAQHvzCnhFoxA0qbeYL0qRJcuK01QLl4g9n1yz8aHUk2+eIsJj
WonLLHTzN51s0NAsIdYQQm+UKoXEGLSqOex6LxDigZLp4y7jNgBYmiRjXYIgncy+pgdHyoeWOhG5
t9okhm0rpx3DvKEClnhrZ7grHz0JmJZwhog0a+eLUJ0ss1GD/6LcxLsiCxCiLDKiabOdCQhLfwkZ
a7um79TBPpb21ZsouJov49GdX1CTW/PftOALHfB+nE8JokNEJTwrER+5G1DUDsdoMS3ZWA8piVZR
H3Uci/Jd+k+TCJX0UonDzmSDT6cJ6nTicZMNwYyYd/c7Jtt33Nh7sg4RNx4qLCwLBgf/Lu2MYAGJ
p2B5VsW/BUP1+XLjdOnqTGH4x8R6V9MloAgTjji/bnp3bwoX99ZqYYye3KU4joVKCia9lgXNZ4sP
nZDySxSbabSZVqavbfnjYSWuKW2dKMk/cuZdOf+yxStt+ZNXLlbwCfjRbloFoucE7l8VFFjuFhE5
GIFhtoVQvzp3sv79c96l6WLR9gn2eZbQygq8vtXJv+YN/ZiHflclVraGdX8NvJB06w0cWxkIOnxD
UaegfvKv7HTkVkzj8JqCY1m/pvE0mZ2loYGLZ4f2jIFXAStOIAxNbQ6IxlYxVWjYtlRy3De8wewV
tAAcCSgdiZTPf2tO6SGgqUd4GmLLDBO4ZIXVYeMuvvkh0Al+mrM5o7sRxt7KZNK2aIQxQP0yCabR
vvAE6j/tjnrTnC/2bpclrDgUAj0xI0TQfuxUd4Dow6fxkAyZs2ZUFoMMX2Hm/xoyDnOTVaipocFI
+G1NlwWrhfIoCFJUrC04n2NRa0CS/j8N0HoqMlmJdzYX3BJ3tVCCUo2+ibJlhw+ugcCJj4ojGrXf
438EdEm50Ikm5pD9lxqKdjr69zp/0CxuDvI9disMgSfvKJj4RwmC1jJhJdzIsne14clV6D95eXTb
beLRMoS5MXbLFr2lLrW2P18pWLcXa6HNxVZYnvtOji3u9y2ezOjdkPt77JW0Bz8+0pSVi+FnG6SK
aNMvU9nRschVzbcVkZqJEbqQ3IqGcphHW4c0FmjOE417Bgx+2uAUDLcN1D3msmOqBzYbV4BHcS3P
nMJd0UDIGK1oJq+Jp1nsvsbvZAGQjllCfhttLjM+Dm7eMhKG6XhF096/9H+6c0CzIag9mijGe3K0
CMd63a3tInoGiRfU3ru+TIENoqoTKTcNWESqA0q79N4nwGy9ebpMSaqr05rbxCW7BZ/1J3xZeAza
2QxtVGvccJmA2fvK2t/g9LmRUddfSpTs9wkyhE3t0IDIo7Ypzxy6t9zHiOwwDIPr2bJfziClKiHw
SXrkJXcUaWwiv177kA+/Oj8S8iVRhmKNfJ45nDK1xPo32gXzP/4hPtGbhc7eovLTQUzUxNayIUz2
QTuNG6fOkzyNYCzvSxBgRTR7NjP5l8OVX8tBadCVR7Zn2ndIDlbuiwpARbPcBWJ3oj+oO9rSiGlr
86U/W0jF9D7eDqcob+iJxJe5HBH7+cBammuffyb5g8JYjG01gPGl+y9iK1QIX7ouSRFgGk1FEC/F
cLfoOlVkSjG1Jb2NOEzSA2/ljgRfLirwIR2VVdT+esjqiKGJoAFaFiiUmZtmmd/1p7JZpS+/g/3W
o57wVJ1ECM/Jxt9+S9gCtmuYNy2BYW7iiCHQHEt9AAYLLjYGlmnCBkGq/2LIotH1Cr6njWcH0+cR
CPpGLVKI68fRvAC667KusLHWcqv8gCu51ut9bKXJ5CjKaURCTZbHL4xogqkMMcNKIOVv753n3ly6
SPM3hnQ5PbyBFOOwTx3rfGIWKJW4Ym47wwxwKa0LvYXCxG+KemVrtaK7cTGrz3hed0tAKkM8unyO
fxYMVbryM0HGJM+dq4HQvBoPdjGQVChCIZM7Fhttc0dct999QpiWdcTWc0p4eIMtvXrhf/TLeo8z
QaDdfL2z2NCjlARaCf58JoQumDzvV1lHJk6u9mVvxZVk9uVLMnV1vXNJlYp/h4WU6oWj8dhMunDt
mKm659/KwFDTWRX7xOU1T0DxoSLuv8d2M43VtTHcBuiUfvMntj/WWSq5BdssUS0NtktcpT5gyxXY
KhYD2SHKuQTZrYFwgt7LUJf4JUcdrexLgwezTY9oex7CtCulvbaRSpUKsm/7T0EEGla1aF3Yvj+O
B1XCXUGxvs5qvoy9y8tVPO8ro6PqiZHa4IaKe++qxS4dQRUa45/YlS12y7flt55dEJPrYYCaIq79
vGn9pA6HzVViaavbN7EW6FE30PBklhK3LBaOZ5Z/x8Lc0pgzfOtr6CH9V7yecKu+Fx/7KSk4M6an
We5dW4sX86EOsJppXHan4T/hVrW31/M3u9jkRHJM5MuWAAKX5FlKmiYUh47h1GI/mmROgW9Zgbve
EDW/S1tFT+kKT4aISb0f0uGh07bDmMVLUpnB7w4NlFCSl85uUurwbi8hWhPq5Ye/1Ql1EyUmZod8
9tQ8lkNPwqVTYVeyX1AS9QbBaJm/Ywjgq01/qDUqFigflygtsC4NcKL1rgzwctnrBaWbPmkPQAZc
msiZJh9YCYdtkt5Akijmjx9VdOAQFBiTb7ud1u19Qh0+G/s9ylHX9YuPFRDXNPyaDVJ0YrO01PGd
N6CpT+zjIzdtHGYw4DEnMDlh1MOWJwD/lECJOCX4ZMxJhWKovxRKGofgSOZz4AH1wX94j+HjfQRM
WT2nmmK+OqlpKybgUNpBJJJBsgAILKsJevprofz8p0XQiDSVFMxKyPmUH73uD90xuXXcUn66Cx2a
ByDZOyFgJjHuE+zveWSDWKzZcXuCntfZY+ap5/ONKa+MATIbLZATZo5GK74ckK+LYHzvy26Sk9el
lYl7naNfYtHCmBprmjKsSqko2xyc/ThO/CWLymy/W+wMDVVwWJOAhaI/ngme5JsDXEEYpF5qeF3q
yUcVOW7+dld4QQu6MtcujHnSMnXVPjwnsudkxihyB/3MVKMGndKNS7lFx/u48aaRPcz7pm6AcuQ8
jJKDx85xQRzXCNcwsdreDy896bPO3DfSfX6zOISLmRVIyhR+RW7kpECDmL7PnSEmhwvrCII+DODL
YOpGA5dj2s1IFGsbgrO6sFh1Putpzbjb61AmQLuSSUKArazNCndfKahtisMa1hUsa0+5R1bklqw/
+VqnDAwNAmPhcVzvUKI4ESoHckE5K9thwBvXCxzwKT9caI73UKLs4AuJFNU1YmEJMCfrWta2Pyat
Zk9SCziOpGrrFYnZoK4tt8I1Yfq2pYvOzgd7Esw69ip+8m4HcstKGTcw432PbcDq4dqRrNVkaOM8
fLeO161rAs5HFp0j8itX9D9e8bykz6eUg6cjxSDHsPTrZY2aOWjhqn0gY0A+YnDv8QN3XA6R2iyU
JvJJ/6+g1EUMo5LXxkBhBbdDusA7NRylj5ZqZYWHVX1ImBRkB20MCAE2r+M+TXpx03z0g3iCpP8g
ctsZuPDVSBNmqCawhP1YPfFVvRuvX4THxKhw8t4aHFHItwFivHtXjimEVtDwE4mRvp4b/aPN6LXB
RTVf0wopPgGLPsqO5yL/iziGvCi69dfZi9BL8Dutpd7dyNlsac81ITIT6X0+frVjbhSgD5ktzyCT
it7dOhGN3nVl3fVAQDd9i66J/It4Fd9uvgMIARYMw088lzlBmfqPwIq/E5uTFLs7m4FZehu8oLM6
v+DqYtxgKbUHufHvpO9q8BlAdjl/pNFB3Gbhz/d7jy05/7b+Fij4TbkiOd/6bogk3NFq4DKdqAS6
vXpCFuzD15dFK+GvFDkIxIgpI80N0yeBbFMVpVHH0+zQOhSvXBbrpcj0juxe3rNQXZpRPOyW+GFa
GwS3diaON0CsXtJGQlfb/0XSy9hWiMHZ7VAWyAt1SODCnYDo/BjZqI4DV4nUs5VGO4sAmU5RbAlq
yWOwH1uxy8qaSxoBzxpWAogHR78pCbMdSpoW0rN1/B13XQHgx8naEN1U2BISSIyeXYEXEuzH8GnC
cZivn4/TQb481hgYMlHOxeWOY854Cjym1ILYFOaZs7eq2tmXXADXrZzq9s/+N/y2t2gZ8dSlmWf6
fI+M47GHfbcvcdwv5wu4JE343M21vfNKtx0RjK4ASXAHAmyZGXZRDL9imVoOXkTLtsYcIFbij3vv
6KOPfhRm+r7I8y0Ufjp8YSZeVN0MwbpgZCatJ1Fd0nW81ede+3FMcDz2z5HHETZ9k4fmgmCgUMg7
9AsLZ5RXv50e85n5zhSLrohYQyoaP8sD3/l5fLVOhrz8brH9q6FWfjsziBr62xV7MT8HAwh6WNIL
qHbfQI2XLRSY5li2qjWnwffolyjExCjIKfruthKP3EjMSNrKhiiD7f3hYzLuCl9c6a/Yh91jcMXR
dMkkYvHqXyg9BZX484YzxgO6URGTqAkUwDyDAe7+yfZl2GBvJDOVfqcTDEeABn/MSDjsviPKpSi6
lcJubnhzariG2tKfeuGgsuLPBYVJMwNR9hIINiy0OeTumE+yqG8UO/x2J75CGKQiDGBk+YJfZ56M
brkxpOINjXRVIu4QdFLfkj8NBVfgB1hCsEGwrUJPTnaq365MVzEHM9wWvPrluvkAJ+jKo3RdyQur
UWeJOe9sU+tLiQyb9H0UVChb306w4DYylXUwMQAdYP/MQnfL3r6uLnoHQPAJHIt3qII35FGGRW+S
oNhvuzJfP/RUY3Zyrs/bRzVyQiqfnb0nE5RDCzgjZybltcRtd+rrq33SpFtk/fswAtb48pvRilUr
vyeTrfTXeF91mrTU6fYjMzFPYfkfftR9vJc0Kod4/Ax7xIyqoywjzhyurwOQoK2S0jWsHXtQvt/q
x7xsSBOPiLIdH8rKVtKBs3oysZWm2/9ELGvIlSi7ljGPIq/OQOIx2cT8F/jTDHuJc4lifjPyNiv6
RPlFvcJ9lE7lWefqMZqcaAtMxrVgO6XTw67ev+USKIVPZgJ/KZmShVI64GtmYW0pu92fqINeWiRZ
XEbX3IP6wwaJ++jQgZ0NX+UFwO6wNOezANomibEcvlq1nYIlH67R7eEwEeBAzF33Sx7MPQGrjjUe
0TN67y41P/VMk8aAYf7gwoGqBk95eT6IZxBqvIoXXAZ35WDri6BiumsbmXqwmOS6lVpObsn+U7rD
z+8jrce+Z2zLS5BLzv0Toc7qXFfEWqTSJ3u30+JxkG2HsJRkRCbQjvqEcNy7NOMxvj9An83TihjA
YsrS9OeqOspyHB4dK2uzk7YPFGJJwkXfaWfQiAYMzaJezQ6yltoMfdp3WJ1V5agjqHcD4F+zFKqd
n3kbMkmNZHUYz/k3UCZYCOij/5joWU6DmvvXTjFqm0/mJMJCUNq8d3AX44eV2yhQyKbj01WNAe83
CfEq3uastLpqlAElti+fRsuFHcgxelMc+lF99Y8RtBQOTeMzmPuBFr1Evoa7UPFFYZOMwSf43x+4
IipFvq9ufInGzc4EbzHyO3iyHFRcRoEcWi3khF21oDU40ANejVaQftIuNJHDU6GhH8yrYISNHg9j
NlnuCk0B8uQxuvuUIalXR84z21z5xgCYyRWimS7C1e9zGwEd3AkN8iJ8sVzBxMfzfgZ5UBVN4azh
UMTqIPxqM5F3HMeFdSquM56++C/74WQJSxuTiEsVu0r+6B6yz3Mx9Wfmb7Adzd8KvEad3A4hSFru
YOaq8Z+W/i35fo7xU8Vs0vNXxEIhrnFsxS2IDRd/Cx8rPdB+fzkwd14SoZHMSs0vpyNVsbUsMW/K
jgAWwesjwxabn6J7LzmAxptxd/BW2hBIcCX9LVvgWib4a7xleaFVzCYLA/PsxsiJFhaRuiSmO4JU
5QIpLu5CB7InMZ95lzvQgABjXGWkaBGxz17W9XuGDU8n0VGYTxqNrfbxsZOZ/3fu0soB/7YqM+zV
8d1bSF7dzvcAxDOR3l4d/N8IL1t6z6qrFNo7CnFskFG7fNi7Al5MYY7JG/IUywUvSDAi5hxAnhD9
h+mv/fBmQe0cKw+BvGPVCFvTZdB6DGq30//FfVNA/z7w9NurdfjDUxR4KWqDjFbTEOocQCXj6He+
PJmiMa32gkwy7YbVBVGqMVR3/C/OvySMfG+GAsyN/gixdEPnYSEQNqf4LJXGEiGwi3iwTu0wfGyL
Ke+b4glL9QfpJmKAQaC5pbtrUhjQjG+1PjDQ0I/bwlKAv6N1tIt3ue8eNbMr93tZUa4qkcpPOe4y
NDwXi2Ql/Yaznlrv+AZB9HKQR7lme4bhM9MV6GiVTxchXh73MvxgBCoailvbOGQ6xzNewpvqWLvf
H6rmNg32R9uDLWgSlyi+KLAVMLnjAVAj8+jDF2Nyh8gXNNuMwSTexNTF3v0zm8tLrLkN1aEZNxrl
PmKECzpU2bwwny5Rxv5gu/UqIMIgx+VHJtw5wpi6MiufkvbgZtumbwoE8Vn1qItGMPxpLNwszgn5
EPaOLxfAXlJxi3BH/0p1EPmz/5gY4QoDc+zYr69SPDoqwAX0wACqjpKlWykmoJirAnm833fTVfX/
lUcQHeMeVpwxISL+jt3mRwL/jIN3ZF9c22DgXUv9MwKH8tKhPvA72GggV/1ZCzVpIxme1dTh1R81
5BSz5VWkUdFG4K6ABKOuwNnRiEr9YmOFzkFXsFRiZ7Z3+n2BQkcVHJ+8Fg4nm5JPN0BqhjpEMO8h
Y5CC7dNETYVjwiaWzl203r2rVCWU7i9qX8f7zIpuFbYTKqz4E5T3MoteiGLo3u3/NDYX7gf7sEv6
PTXXVIspuNA15IgjqJKtNCqDG6DVEuSuRLge9GBrnW9+Fy14LElI0HsELtEMqotKNqdeyJ39aUoC
lCxcd+kti67ShEnUl7ZCyvOpf7c1aaXdlqvgKB6LXcYD5L6EZKdL31xRkGBDXHDKlh8V4ZLiHctA
DH3kCITWqtwBSErNu+jDxuXALXd7LSv2/8M0a5xhSC26X8d3bXj6LXM9kICbfhEf0WwNt1AaK4b2
S1EoNW4MBp3nUIoa8TQji1C0+WO4DHb5DYQqj2Rcm2egYMWO8F0HsQHUNusoWE+49jM0/2ajqLmu
HONOOGSRaCstmJ5QwTeaQ1nR7EhzoB8F8XcSpDZOyrLBbxauGoBYFZD2BJrVadsdl2MJNdApLbxZ
dVadjECsInb/3s77U8axre07q95IXb0D2grtBIK6Fg0nYchQ3ceqV/8w9iLFWK1mH1Fh9gk6ZrXi
LDJood5uqhkoId76SnGlXzIfMOfqTYt3YUUakpraNBkiSaGgz5A+A/CQqCI0DCMS5kmOyAn9LN3+
EHMLtZ9m08ze6PPycoQl82dCdC87leNM3LO5jAmLP6glzi2yHZ9GeMcUrTmA/6TKHDt25VuTCxMF
7en9zrCYdHlLWdIcOc+ATIQHU4Bn/mywt1L06AkVDTqTA+/PLA/jfiaSRBI6H2ok8DRmFyAENrNx
3koUfOE7Rt/wKNoMPJQ6yDS77Swvf//1EWsmVVQ98g4eZOzFLTUbf4nI72NLVYHWQkVVI6rgxXH0
7ajjqn2xcfbmMLEoAQpHYIYDZVr1+9Dk50NtBFkUP0ZZMYwxSqOQoTNwvXRJR/wXQQKSIq8lhjWL
uuYnd4IW0wuh6iwZL1czQeCL0m5IbwDIgvFY7Kl7HfQ4hXwbw76e5mhvd4xaYtBRJRuBLQWx/Ba3
l4gX04ErXZpzqq9n2Lz8i2zIVAP2lmqgI1HhpiKv1oBAb+CDJZArqLo0BIQ87+kiTIwJ4NsbwYUJ
zXCHQ/gpwFirAsYYrGuHJ5KRAfaEX98jU6IJNA3rz3VUw+Yk7a5XBD6K/S8AVaWKZ24zFxI/VOcu
75a0wIcENOXF1q0LV+wjxHnTAWKYI8FHgg8q6HDhNqdDmP0gblKk1E0vNOwQuXY8XE0nGW+kZyQJ
R7CpizYPWmzgPbqGvjuAA0PC7f5qPWxkf2zF6rR1sLNLW2MYxYV2ANFoNHM3/fUv/f4+WDW+FHZn
/ltISoWMLj3ax20I9ypys92fUck+JEPIlDNyOkGojZK4vXP4T4fo/GS91RkvTz6qG9mK3MGSf+Th
fR94B2zTtrzhjR17tq6dBgbQbrZaZWnWwyX9p3hXae9eRcHS6N0XYFa/a5Kt3IvrYR48lh8M0DzL
LelccS6sAV33Z0TIiFTvxFVzVJEU5jZh4MaM45Kio4TUFJdf/wuK6YaVjZsHvkc3QYzwvjWIFvVe
s6p3qsi48EB4nhegCzR7fy5Gys56yrHT4e31B21PGkilX9GB8q3mdryH4NALrRJGKPXBuEcPpbPQ
RC1+g+0zO/mTnFA35mRxtw12UNEf9SrL4TCDLQ5ZLzji4TAqvFLHph5IFVhwndMHPvjYX/Duuhdi
HbsVv3ly5Qf0SC7fU1lYW3WsEm2teq+IV/kDpabuq6LBABvx0VJ0jKd6TTSn5O732PJRrk0GNM9L
tEyZhcfNJ1tNAgGDQ8KnjzH0n4c4wbV+vGhfbNuEScrzAUhZ3E35wWjvEqxAdmclDIvYyk1un3lF
gGY/+rJwUAFDU2M+sm3yDJnvCtQpIYI0JsWEuft4LCvbyjLU9phUCE3BUvRUfhaa4shes9AkWKm8
Rw0E04F+I5oFgw7VOQsWOY0McZkEKm8qiNQjejWUybyiTZ0ik227iLg/Pw4caDGxgQ/tFsf3wnTe
Js+ApUEh67zenWic9xnkGtiCJay4zPhv/x9+fpbQLDGSEDUCEXpCBH3zW/dNIP6McJO0yI7QaYn9
IMIeDv3yLLNrFm+vg0boQcV+Xjb54HdgS4zioVt8N5tIOdDlA0K7SrpXiAjuF8L4k2GWCwxTUVdX
NY0QCJUznYIgphKTja2IOiJH8eAvO6++NY8QWI2RIYUKlBC7+w5RRCIbQao+Csr7FzyafnjywbKn
d1x8tvcWqvQ639hv1ikd/HWkjwIJM3Izp1pvVVS8x+ZoGH++cqS4VP0U/hpGFjXUK7QHJAJH+J7L
a54DqAmSNCMZrfCBPJSa7UhJEZEsKjQfjKbXxbsvo14OnW063l30kig22Tz9/VsPEDVe432F01KZ
hUQTjdRgAusp0YSrO1oN/AtNgTLcn4lKyXB5E9JXL8DzK9pH7Y8oc7BuIYicnZmEduVS4Tr1GWNf
paSroxhgBs10eF3sJKgyJDQ8f6iI+6uuxt+9flgV/BV5houXXzveiVDS6ZK6aVnEennDZHX9Wo6X
gVhqvlqVNkV9meWBfAGlna3gHScI1Vz5k/JQ3E5U3BS8XeCzF0pQBl+zgag/KdD9fkR8u8tsStov
czK8/O42JdRRVJHUtInVHYkOm0pBM/IDrHSWOhwbYMXYv15X8zRPVsMPtHaqEcL/BjSeUlHK2tIq
yJWSmiGKLKl2DXyQV14q8MvKbbUxEUZNH4nLW8pHMHWDc4pnk4zwaiDfbWcFlk2GKPpeKEDkqNmI
2AZ1X/hD3eVOITpLIBUfPy1OjqkZ5LeK5D3ERVQFR02XYxu5gCV4dtQBL/lZ3mly2wqErcCTmCC5
lQ5W9/l655G8cTiIPFTcR/8Iit/7aBEPpQTYzhU2xCGzmHL7ANyCbSV1KM2ibGpIImzibc0Ea5Tj
pn+NJ1h4U952iKkxTG34INzaW9eEnCyO+xDTZ2ZER29TSK7SSfMbj6NyrnRLnNm8mIAWIAw+Z7ro
iWgJG6DJTx85lnBPMsrstGs4O5/TiWmAD7jsL7Y+7NXWAlFld/knU9fJKybcucTs4N3QsdwdICq6
pGGvsQeLZHzm2e5xcQ00g6//vq8he05lBjQMW3AhZDMdWjDkZM6OCYar7HqcNtAKu38vwPDYxtUT
gAopmB63UXXgqGSd96ktTPdtBAfJF6DAKsJRYZv/naKaa0CB9EOevbTkvc8UC/uZNhzEIbFKWOjr
1PKpnJA+hwxLnF51E6CHTpVbhh9Xc529lI+x++h7tahKQeRumhR9VmxETOA7LgBzq1xuzFmCVxiB
hSjssXPOobgAObfKFVlNRNfJujpbHgFrWVQuYbMEk/5vwGl5komK29nAIKZj86skQQtMWQiSbgwW
SoVq2XJYpQE8pq/QjL2yvJxETxS8SQTMnLZBVKxICnPp5eTKpsl2XapZbLEVx99R4lVV3PEznP9h
Ae1jb1vubAMwU9D87S6J/F5YKZg97WewJYzcxtNfBx5TUUOmV5RmXgFUoSLgMVxqGbXgrRduITKp
S/WQozzT2dTa2WCk86oELnFdrvQggB90d4qHSz1XswOq7z/TyXKqkN0E7FEaiBBKYd84xUKwUHEv
3oSO+AVfIfkKRgfuyeMznukd7QZOS3SB6KaFplMI4snv1Vcgic6uGkQfX4kVtEL079dJwwvK5jcP
Pw8mdH6VawnQRVqWamc050ymcBpyq3clAnd52SxzgXoAUch23J+n8Uf53rhUx63JhQ78TbWou9MV
auSlLia3UiE9O0km3GFoySX1e0kSJSYh8dOtytD7F82j3g7U7jc7ANsypx5qy46CNoz2E+QPXObB
tm6aV34NP7kBjs93WwLh+yeq99408eYFVJmSwvxOIWS/M4gOG+VrfwbUKbKO/XLyDqjb4FirAdHs
sfRV79uHRUlW6Rj1fbx9Cn2HC/BpwtplzXyROW88iP88z5bdhMXeK2323XTT+zqvdzweOLzgnZf5
nI7Hi5xNN97dB6WsYfPVgnkf+oLto32/DE0PgISh202LG3iH0cb744yLJiYsh4v9HrBYJJ6tVDze
XMjzKRG6R2/KK4kezEbKbvowVsro4CRQblKX6PqZlIjTk+ecsfqrjwv06tCMS7XS0ce0vTxQ03Qg
zOEwsaFwcmdyiqHCs4Jj0GmNfbpMFyzasppuSaohKZMbSilcIuAZEaoDiqbuj+msTriutEOwrPIU
G/j0jPZOKlrEV935eT+1ts8/F1ZjOhoho6IYZL/ij7QWYL/rccDgiwwI9KkULL4BstebLrKk7E9d
1c2IR/QZEWhJAfXRcNYBaOnMH7Rugy7cpuAkgwEhDafLyYsqOsQ/ES3WbpkZEbBQvWRxJQRAetST
aRbsW1ao0VlRKpBhT+T4Nt7Ltg6ZuGRjhBYycAxSdwwtTMwxj8reqCH7p4FkjowBquNec4qCOCF6
YMSDkFIRv8gUCmHRlAGhFfEBaGV4UWROQyfh7B7wEHLtSXrkzIfhiY6ItAmiYlswEbOa4KYFzrEc
B01LaFctsZV7OiC0JPasWAh9iOLJuN5hEG04D1LVyoUtbkqgJxKvKO+En1i0mFEoLHGZBWk2d55S
IbdSVApdmzaI7ukf6e4ZDaFuM0PCCgeh4gW467PwZ5LYZ8RonfwkIptJXewKpEhBfiISrK3MuID0
HeFGt1Zv+yrTv67REyRH507XpEFcBkPqq+N+BBUCHBHdF7hxyTSP787e6WJE70wyKNgaDbdu5bAz
XImxM/4crQXXSnD3VjDDsyeqeUy5INyhlQWvE230QsP6LHOhDHDnccuo2pl+06xRCtjJs9+X9xCy
71OPXUvyvWC2HVFKAtUlk6iXmgO2bJE0/yzn5Zo4Y3V1bZXO7jDoCewGVQpm0ZB2T8u3Oszo5yYf
DI5ES+bc2vD07v9ET855btT9CImanEUJqoMG6VFWVNQ2m6VDp+ulkDK4CTjrKGrROQh2RIhpbOLj
f2xxIXDLGX92OH3dhGu5UpkPYEbxKW/lyh5c1R1iCjQxhbeAoYwDPkWED8ZePygsJbU35ibkx9JM
cbqnw85BI/ExYY+iQKP3r+FZSBGW5zbGGcGPOvbAPh0AkM3HM+n/D6G183Xrr3oLeqUqzt8YUjbW
lyh3XRiylxDRuWPtvsH2dxaEtLE7We1irDmOBQqGbT+qffk8fI7SXElhj0g1E3YqKYVt0Ffw+VoG
gecivGwnFPzDNPlpNXds6Swaz704inH+2BF7tmtRpprGoY30m+IeJ1lBttLzVHCt6nYX518If18Q
ZtQw6mjWmX0mB7JRwBAEB4vODf/FOPjnU9bOhxE7Ix1w4vODk3Aleqs/0JcS/VckBN3xz0mfRa64
PzdseuykH+XmZBkEzFUC1hqKSnlpSVDY2ejTGb/eEch/zFdJzRvg7NwEEg4thAHuVfMzRzgWRoFb
Tk4o1Eo9WBiSw/fd1aWHLel92tL1KXIhZVOrMc+h4pDzCYADJY7fpNt9jmqFuRh37/NnzDESti95
YC8PvJif2vJq16NvDj9npOZ4uTYApfVXssdPNKlzNz6HkbNg4Kdw5OrLY6O2dVgFkFAqj1NqpzVY
glXtSx3EId3DsdhzZXmR6mlgwYz8nbJQUMEPMP5VZom5QskWgGD8Z4kkW3kZmFJCKUZBCujGErUl
jGFTK6fODWWYgZKUvvUFKr9mBX67YQcbUQxD79NPPW8sAL1oypNSO6cxA9SbxY3MdR/zGZBcgNGm
dCaFoH0y0Ua5HzpQhGIOS/iFNgrD1Px+ewzSBK+vRyYKOlUAosqYCRKkGZiinWGJA5q5FgJOXf6J
R/26x0KZiN4s+VHQA2D3oUgv9UC+yikJa2Z2i5Jg20BGrJt+Lnc/+V1yH5SKbVC+YtvNmpn4+KVu
3TEdH7KRlXBDWh4jY4f2AiRugOjPA37f8yhCMR4kFNf0U4bId2F/fCWQ30e2ATzxtOvmHL86Zi+3
N32Saj7/3/FFqb/rEWGvLTp0m355Sgry6lrvuEzyf+xYpqrXpFpChulIVbFblQw9nnpqndXZQNWR
A9SCobPRkAn3WPCSL6WWxZ/iGvk+SXhsNdpAqUbJkuFNXIoEAVDuBk9/qRRrpsPbdozp+cFPDzgX
1mN8HWWGYmneEqd3NFqVMYJM4sFHf35KUdae1o235VObT1p+WXC6XWZn3pFwmjva2K0UI+UMRDXQ
cpjJmg+jab7Ve4AGLKntVdgqnk3n9LRtWzzTWwASbSV+67Buyf6oOC4nzyEVtTw0AaVvsHNxRMrq
9mDrijvPZWbWh0W9k/USSUDJr/6wgGZpZ872Pk3opvX+rdMwYSUf9PoejysbbSrp6QFnhtkeo716
okakD0Q5b4Hd/3Fhr6/7uo4wou3a0RgEFd1od+V2xrOf8mA+cBOR9Q8dNz97MFdR7prkWJt32R2Y
2gG/sYtTjzLq919+4+2aJqfsUp9BiFrg4JDaZ4OAJfuKE8j/y6NeOqTDgPfYfDy2jrNeHKlXOmT+
OkVM6VwjqWJN7hSECLq2EQKFaAcLTuqaQY0Mx+8bwEnhb9vAFcltTha9uQI5hSkq2bXRDYXLkr1I
+0PwnFW3J9BRqskysYUFrGhr/hTTToyuXeU/st6y1HGo0W3Ct9ZSXijNrpuqXvqaz91rSUfFKsgC
DJKsrA8bTIL5m6mdtBkKo2a+IZhzGRMFIkDl9DBQur0O8yAmlY/SexLZgG8GbkRZ4I6NYczPqtiD
nBOg2Jw3Oz2/f4cUBpgge0hrKQDKV9l96nvLxL1h628WyMqF5IFws5aS4rMBsuS7DILk99iPjquq
s4FRjzrPSYM5pjGC/VYvKgdoDvuSrW2hUFwQa9vUYx6pHLGB7zF/YB8D4fLqFQI4h0PpTgMBErLP
G0jbQgckNwPmvN4jwgcBlVHXgT2OBe7UUgPRZ1zUrAe8L9MWsStOsxxe0VO4e5/ANl7CQIrNfwZn
/MI30DKHnYtfRFWCokmxRejoHXflUrwWg4TBJ8KshlVreSQXo9SawYMuqGG6SXVictREiBrrBIIg
bTtEs3sn7BSfPvy9BVhFz3rcBOGM4hsP6CsFS9Dbm4zs+hHEVS9I0/T94ObnJY783GE/apt/SCtV
xi1tmGbDF0NvyoPuw7fbD/DJJRbn4Cro3qVs5PKYmC3Zz5vxEBAgwDWOxBG0sAi14R2qvBQrh4nk
O21zymuhWXlq2fshgjOoNPDUS8TbU5AdhLHbT0aPwH84ZEX44mjOUXUvnruDFxe8bRl5kkHRmguu
yFqkpFNsDd61vlWeJDdI0krBUzhjzODV5AJx5B1l9xmgTD1UtJXQtPdKmG8RtBWzQiNedSva7xin
b5uddw5uhxTwFrTo8P3LtaiDWsVjsTjRVVkvmzGd3lBjlr/CWuLMCPXsaf9Y414YJc0GxKbHYdoU
JrFm0PoqMCIyk1OhNUEHb1AVEqjPcXNHuYsC1kDtw05ZKIDG98LTHxgFSu6hHVw3J8KUHh17nm9A
8wsGeylzxCzusIP8XOlF0qjf7bPVOCpHjPIUJRDepGRrjJKaAG65n4SiYU0MbWZeM3XSG5HHQXfC
NMHTGgb7AfeVApd1MpDyU9k0J/txFLaA05PjEurhvDSrW3BnoXsWUvMZ+N0fY7mvlg8BMBfkNg8Q
i4VDNZkHV3RpuholyYN4Hh3ZpV8emaLcUNfG1gdlKdKLhU5IvyDxoSCueLOABrghLleoE94GDCwH
xp5UW05eksv8ARnlNs6BFFgfQgzXR7NERR+eTp46dDBgVzuNTPPw2Ue6F31OXP5WrCkrzxsP9KDc
ZBTADf3adzn5MpGpI8dL+JMG1Ty/G0R0P3PoMo3rUX36GpfOjufY4LgxkdNyx7zewVeNGqFuAdL6
h3x+ycoQUrtwKF7VRjU6jMZIhtDisMOC0mYXduv96EpC5YkWxsOpFVHYB8d7Y+Z8fpA5T6FcR+L8
RgawvYXp/Rhxw2iSBMWK5YW29FFWGvG6Ny55Axm7Kxob8rgdoRtm5y3wp6wsaj3UgKKvEBhmYAPz
sPq56WmjP88KmwvsPEMUevufLT2p2vRhicWQfdf0I7ZB6tgJYpVaQgmN2WWvpw+tpZmhc81FmiR8
+e7q2AtvvOR3LqPuB/nV+uGc+wHZ8lRoeVsEkeIdJsQFlCJf6NvinWczHDnXeqOXPBVdo9HfPAeH
+A4A9fw1F9NFk/X8K+ivaCnSMShadEIBjqVnL1lsTOaWBKareOJ9W+uBOVldjbg2cedLDjPk3ss5
LCC7LuEUxvaes+6KcCyQJqI1KAzee4Bu9v7NsKOUyK+6bZYgqQJ2fHfhWDUBDlzrtP+2ceDT2Fbv
mtqRLZN+eb/xNJftG3GYnjkr/Np59ogu+PaXXMa8hpkMarXfyFjH2T6zEBrQV8bkrwphE6k+BoG6
D0OiXURIA6/2dTeaQvGHWqE+pD5wkk7KTAlWTh8QyI9M0BltrxR4h6janK2/LH7dUK2jzSL1rNus
d6UPi7A01NFIrYJPHsLH1GuuviDCS6++BGXVz85fw+kCK/RsSimqOvEE+mDc2u/6Moo9sGg6ij3+
B0Ikm6e41pxM4JrR76MCNYzFkoaw2kMmkz8H4iXCNZgaWoBaLg3nyzrwqsLfbVZCOC6dtzhXXPHI
5pJBtcQG+2sVPc0FjKcr3+zGlOhH7PL6Enu5nqeIXkYHSOVwJYbrXFpUZEpty/W4K34UyfZRIaDg
GK/cXiYU8BBsHCzKnp8tm/KS5JF5gi4obcHRHx1yWNn0dFxW9YRraaIstZN55rFbCj6ZzauN3LYR
Ns0OHfrTnASuqBBXMs9IJdyzI0A9HaCiuCGjCEEIt1JoFGU6utaEmiHsqbVFr2BmLQZJxSK8fhpg
tI3DXzwz/WxgW6Fr/T++VSnitEmmqHNOQLSY/SfPVTT5sW2S8xxft77ttjRgJI+gjx3gSkqr/bdJ
GZNjfyf73oPUqy+1mT/9SatEJk3q5MCw+fozwkL3r3j7bsf3Ft3Z+bWcbtOGgCj2S+RqGqHWxuFO
FS18ymD4yv4NAOfSeTkhPmKDyDPf+eEXiwQdZ32MZIwy/0MIr1esZc+H3txpPLHWqi41ZmmLeDQc
C+ApnZzyThqmMEnnOHppn4lgEIyCiB/uKwDCHm5w216zEN9A+o/ZfAZvF0LI029tGpnwREX4MjhW
iaJ3j/70D5cibrJJabDf9nNwdGtjHLMHHqkAd9Na0xa1QpW+sNmuXE9p77cdHwov0KHjMIOzMvWo
wm4yhN3q+FINZXuQAre07frYMiJnVi1tHaPqIht4GiyZcYjcJg4yWhzg+L2ICG8VcFM/vv5xToYh
9/PhTZUpvfeleak5dmE5x9Wcdok1fk4GRlRs4MEHRCE0JHPtDpO28KiLFVQIknP2hsVIVueMFfom
rwC8LxWF+Mhkr+tKFDCWancH4EUO17G5l2dJLTWGCPA2dPRC/iixc+bNVjiTDgAU252pmv+sUoxB
00R/hq5psLwL339fP0nSi0QgaqmnOr45bAVytCD5s8Oq5evYpW0Zuj5FAt6LOAeyoJYo4OJfm2tu
T2xSTP+S5MehF/7Am+1Fb8ntbtebnWMnhzEd2WjfkF4YBata9rsODIeBXfr6KjfzcOmvR8nPgGvA
FRDlCr/ANS0Nv2+sqiL/dHLA+zLliJnAl0hhxgX8OJ82Xkd4zM4+dxvh06FOjfu8tBsVjdAfuH2q
Tr6mcTnyekBm8v9+34z9+TXYjXR7qfM9QK9GzF2rgJ/crkU60Xh/a+6+DoFWtOAdsxfK3JpG35xW
hFkEL4cbh3NgKEBcjlnbsqWSa/5KLXsqdbFeF3gWw5+MlciwDCFkdFg0qQtcVAcucXYuVtnEyWj0
ga4cAJvISlU0xli+dSKX4r74k6PNIuxata9DYQ2k3iHSUPT/5CC9e3kfEY14kbavGgFv+ZbPRci+
0W7s4apwIASjd/ZIg/7GbN+U/JGf7ttFzs9apAD+YGv7U8MFWl/HCh02USPjJbdW6mggQ0qayI1k
g9brv+0xl8tEl55PEP6oxjjEoXHe4a+C3C8X/H5vqLHhIiMw0kQncZB8yT3sMhvlo7pClKNU38zU
QnnDgise3wkAHA6R7PyncSyUXCkokcikedYYJ7kVOLXNNSsfDf9c6pKS9Wi8yEIGRvTtWqoXoZO4
4iyH6U6p5A7+viHN7lXb/+V8StR1R6kKJrac/bAjBP9dGHKJzuQh4l27wKD137DJBJAA0WJ8NQAK
UHduPM6ING810Xf7bRqiq3HlBJ4RdX5Dd/WGu1VS7dSaXhjgvOLn5X6tCOX1iC1XhtK+aSvi4At8
2fEkPWRLNcOwcVj2jOObh5lPMhQGQiTqb04fWbYzjRquBl9pYTlMQfJoVbKpCR5dqT+WLeYSNmKO
z7DN745gT9/XamL2lCSaV2oDAG2TMcqcahd+Po6NyZ3ZF3X3K0Hdilx8ZOjJTsc4NkMNgoDv6cXi
PmkhLl9c3c8+BprZwjukPPh5zudJ6t3G5BTedEX41eyMF8CdK1w4Yqz52DS9P+xJ4WAgmt2XDsR9
zkefq8Q1JBaYOoFyhvmb6fy/8wH6gMxPson50fs1riTO33TQgnGplqFepJTffsaqwjthz1t54U5u
05CtaVU7bzhdzbZEhbsfh3DdEiqDqrK0qIhPh2MFOh5SCZp+Cg7dmpUiGwIdLLblplQKy1TrQBG4
372uLHkCMrsbBAUGov+1bHXSY3cCkJVLaoSNs79+2kMZS8b7XrlGHaJPHkmKASnU6jTKXEjnmxVR
OpBAvcHXom6lwiDs0+UXpa0Dl4py2R8miprkil1zrCx3DhxP7X4g8thFUuHTqzW+WZPAd0WoPnSp
/NZLKcunl9vEfI7jov7XH5GGTerMDx3a6l/DxhHVeHbieib8F4FNWf5kX4vhh4n+QQyUGiFsfWWm
S3vUJSrSLyiP9QKUhVpaCL9jQ4Wu9OGKbfd6rnI6+SOPRMYuOpJC6qAF005PKX2X2FjAoxamouGB
YXCKxbu6r0IRvcIUCt1JTta1NrkshHnwqO6x+vxxfIVoHooChqLZGd74d7quWb+Bd6clofu+M/tI
dVZnqBgIAt8vbtNGROhFif+JQjvbioDhwVyHYK/lA0d+H9jYdWpeRep5fwbTXssJo0SQ2MtBlEp4
atsfKqZUynBjwaBJw6pG2ePdvUgpzVByoylMMJjvk4dAbHF9S+zG/qRGubbdVcvGiCU0BMHu/OtV
SLZUduW4bqHddlfVvoQctmqtKedjCbYJjA5HC5o8bfgqELRoN8EZ5/dsGjHacGGx1G6eBKsEI5C/
58QRb90bpQgiw6XEsFGZiDaMb+YAemDZd459Z3/D+5VHMZVedvCNHUw9aPpiuZdXF5tFanqRFahC
7TufroKrckaZ9nMaYcAvexrMQz5OrygGIkJdkwb17bPKPdQw+61w4235bQ0yRtjYAeaFXpLG11J5
dq87E6VttoN1FmSzd0N26V5P0GuuZ0IaJtX3z9iYdGGRNRNOWW56iyY4yl1yWDx1H7kc/Ju736WD
Imnxepm1YTA5DDhLU2vAhvrk/Ke2Y3tHj8SAovm91nJhP7GcOgyLe5++zTdgKFoZX7YDPSP+OkA2
3mFQYaYUlC4NvzkMfJRmT5Wo2l17YHu1jLk93lyGcYbiyORyKQOd2+p+cY/APrGQVbM71voX5TYn
l3yKwxuALa7tkRecFAbv4HFFuDRUKhQE/JXekC6udA16u7km28D2WbxSUHZznzeCuhub8tJZoUJb
l2lbHuJD1SDojSHFJaummgUqH+2iJ/j3r2+j0hd7mHh4qyu7W9X183W9wELXUv3m//mHIZhKfSmb
TuFyvro7yFDp9aaXYplzFbW+yqJ1KoGbyNGmZ+xg7VcjGCmwVDrmppx1w7AgfKI4mhf4hc4dZ6AC
1ySpMW8q+TS2iz6ABXrCwW8lY7P8lqywNVFpPdfmqwJaAIWC0zs2DKwveFOkqxNbfviZGWwWTxzw
u2Bo2GOCvafDvt8xUJCjjd0Vu7GeV9GwT2Zoz09MMXjw6icKSto4a7uEGHEQOAswZXU7viqbHVXv
C2J0N5i8b5GyrRIA1/KAVQc/jOHy68CkM7MVXospuSTujiBsUgpUIr41mQoCufgHqKVJOw6N3y9L
x2jl1K88RYzumT1AOCeRxPw1Qy6WYkkBsce4BsUPUxfGRD1L8C3+lPe0nXFMohNQKqYNMyKRN0Fe
/GFPR2Q4+WonBPGYZvI+fYvfTltLZ0I+QqfRBZtn/ezZBjptAsdBOHmNJL+3WdZ8idIZ9TnlHnSM
ZCAiQKWhDscPexaMfUajv7sVS+zav4KdZsoRYW6ZRduLakPL8hP+HDj6QwtNAzydkDILgGaSu/7a
GaJhBfOVjwPpBJmBam43OGVKDLCjKUt8lUvq/u0MRANwg0Xq0i86iCkl6qlC+uVUZPdi7es1CfGy
Ny/SQ/pIG/Zdkj74lm4fPRTmAdbJrFe5JtUq+bCq/woCIOuCHPgsMnIsG1W956sryYqRKXDd2bTv
9krjF8Jzba7dNpZWGAC6dP3iaA3IbNUM+dnPhCSM8Z2KkgDmlKIrqi0GTR3iD2V1OQ1GnAO8NHw1
DCIeX1u3G0jA9LLKwmTwhrBDtMxWpb3CgDLO+gtTgj3uCmAT2mn3bB/vynrwTT0VRxtUn14ooCts
dKNB2HUbryHte1rSCSPW/BmhM0DHAkyeBZghgD+QyzPm8fOC0mrh3m7Nt/ygi1ltNuK1IR70+N/g
ZECjSxskoAGfVLaxp46AfgQAd8AsPoO5Q8V76DZK9vDoFkHMijTG04RjlHWiUA7QuRmggiWqYPAu
GsYfqY8C/olS2dB+oJEpPrTpuQJr4H5YqMM1hFAu+CBX/dgAMzRjjd4m4sTZ0iMfL8TdgnrQXLjS
DOy2QpO+the4p9de6FLfrlNtL3as8EHQOpp/zIMxLJJoBhkm7pIAoIgR7hXDz4zYQZylTIQd+3Py
9jhFfNgyUTahMBnRAIJUBQX2Pp8i2FvzdNTk7HmFb7d5m98RULbsTs4YmKOYzwY+fs8zm899gO/z
Bf9GIRFG+A4DgCrHxiyM1Wx1rFalG+E9habLH3LEDM1x3u3CgSzBGpyDbj+rx2nb1ACN0oXK9aIP
5Pp/iCNC1e05wOKkf/Ed3e7Bl1qBmN2wiTBsa8tZUE7uZhH2L2RfJ9onhZIq8dYDw9fwbqAbHEeq
ApWse9pz7DUvswlu9UnCmRH+4PeOQIEUgW9L50IO6sUlpEkRfpmILad0FPJxwgvG9sJ6pocWBOR+
kgVL9dTsjV919th1K85PNBL1fZ82gEN4uEguk5wQWJP+KDkD4MEo5IVyvHcnOHhILY8HvXwQCYeX
4rGp0hzTKagDfJH330BFDZDuL30Emo8NnZ5w35mvAKZCCAojCPCxY2AmC1FzT0QrVKI1WpVtM8Bn
v6mIr+WClWMn+nux3y8+Uq0Z5w/LLT/u+wN0fNbZLMDm0rnX+oFENUJDHpvWU0E7/U+CvJT26IQd
B8nFP/iElWkE72fkjmjBpfibGCUxCZ1b+bvkiOW+TTg4SuVbXaKNbhX6h6n1UJ70vJVylmwYjlA9
Zhr8YE0jbCStysc5vRC/SBK9MrbE9zAWJaQZODqrzaN89Li4bo4XHf9HBY+CQosn0cPZyswfM8tf
sGIt58ujBK7e+nDl1t70mOjluWrcwyHbvJ5z3wo3Jw33VvfPjtdw8+KqaiMhiHJGKm2BewGBaYBF
bBkNYocn1rOkSAdenlKWRBsrtkS6NTTZcWepJjdxzGPUI+8RZ2hSmIyj3RVk4xLJdgV89guk9Fto
k/EaWeP7qG+V5xt+YhmreNPjc7ltcsitJg16l+Ux6cCo8Td+ljj0EW9aypHtZ3qqSEb9u9OOD6/9
1C94n9crg/RobmZWbapECkXMD/wuQrD1nKmKHMYf3NalVQwOzENSJigXaAvOl8p6tXfQpP/qNOHO
pzNdRphPBkWwjUHN5hsHqumo42yDes9+Grl88O7WavGQHy//vv/OgkGZNKtwOiB8w1UqJVRAlwoE
Q+CxUnUKDztOgUAp/K2bNr+nVfS5JlYIRbOiiNaMKN5+T3xs6bpr7jpdLh06lUzgCATyWlcdBsWL
Dg0Plp0UhewpRda8JhLNCAOG470gB1dkY2vQqJhNkZ5CIvDeMv4hD/6hzQMr2jLVSmRqJym7xRu5
mynwkLuGzlZ41lW9UQYvFDskXKA4ytapQiLJPhoMfZtu8M9TmhpQl69r2xy3nwvxlEI6s3+3B1tU
BXPa4mliK/hSgztC1+l4hVbPib0GB96vmJ1erKPleEsuMajbyAWq/VCBaD/5x+6FUaQPidz7PWJy
NmHhP+YO1lpLH4pzmx/1rlsibk9EDhD8E6rK0QRnN6RvVz/wu0U66CRrGnB3a+GRsFZhU4+wNLtu
H0uH/lHe8FDF9xpsbAfFl05adev6KcfQADvDi68hL5STru69pxtr3Fru1aYwd3Oefj7yHrFm1qTm
xgWnRdVeiIzKxvcD+VmEFCHENHiAd1THDQDMEyL0QaGSHPVIP25dG4iO2BINKkqGQ27OAkoihATF
+F14cpRA8zzju9hmITloAwSMI5XJ3cdkodA3S/8x0PatAAVJQIf/JV5+4dxzc3JRWGAhyVTkRxzf
xbhEPt3Z99NNOfk25MDjHZfYD4njCCmB9tv5iVIa+8uix6v9pGyosGg5URu/sjmooDyzvGSAxHPY
t6/IrVZ/nSeP1b+5/5sLfwQQ0x5cxSh2lgG+bBdzKWohM781sRL2JB5MfM329vhlNRKwXIj9mGlk
xTbhi4kU4+C/OQwDV2zOjZK0xs7JB3qObaO1BY2RUzHoggcSt71UZZffT//ajATAXiUYvR5GMl0Z
6qz1IpREOqByHPJiemedWKNG72H958eCKVklOYYH6pWI1nLe1QzXA240Ww/2QJ+gmR+6TlbwAue1
Pl3nTZjuW5MQfyp4Vy/tJwQH81Xw/bY6/xc3qcOFVfevjWFl+w1safqTVLbx4N71bWbHOnt7yHm4
PBzGrYE0CQgcAM1lKZzanl1J7s/mHIWweZcFEY20ExPt+8StbGsfQotpO88bKtBxClXzlHdNjjqV
eIdIBK8Q14dL6fnXcQZsf8w5QF9bRblRaMWtqwDcxJoXGZBuYyBMSm89tadA73jMyFeCsU74D/pv
7hND/KqY5AOPq8EAqhXVCE8Ye4y44qyi8Ge2jwhn/ah6WjQr+C/I5aXGHXJ+fsvN67dNnx/YhxVp
YSbQaUmaIhSRvgxM7clrSdOJzXJ+POWfb9EIrE1K1Y4mXfJFGaZRlH2tO7oE/SqMlpty7DPoyfZh
gOqmxt7qzgYOYYGYhqmLlP5YbUJOsvNvxaQhNdj56dpAntlP+Hc6it60mGZukMILvaPj2gT63iI/
paTVkIedQkWbCXjWPmr5UaCHsJ+FNIRSx/An5obWsOeGQFn9zIfDiUR4+mYPwLKLZ3juVSwLgd7Z
3S82/RJ2U0xkJxrqYCtyJMJal5ysH/RvBbTgSjnviuwoOdpCMO5wbEpaRCZorp62lyhynmPdhO23
g6DN+tyfJwDpF+XgGM+8hJ4gJphPG1k0NMtjnDzzYpy4qUjB+9dEayHaMOIQp2bVaXkFSON1nIuL
lyO/572sxqXp3hg901LnF6mFzCviouvHBKLJYmjP2a9FpCkY6Xoy2bW4bTkeSVodead+vH/g+X7a
cgo2bbIEh7GA5IiYIIQQQ0laQJuG5yPGu5jjYRa1klk7/G7GZUDe5ZTjIzKEe9Q/GhrXAbmKjZuK
JdKwTdjgIqrdRSSDt4KtjTmstaFa5Sgp3bDUqa6feLeeNTmfoE7A0leu9SkXYYLu8K96euK/P7Mq
SjZyDMHqGpUn2JXwrTV/MOZNT7crM0Ira4YfnHRYao2ekT63U+Pfdaa9Q9Boit3XberMRaP9uoUc
kEg2Konxdgy9FHxzDUqSRn4BsEp3xfyK2loMMtd1pICUcV6V2muWcB/ENxHEcToOC5cGzD/zNw6/
8w8hfMmyoRTjKIPc6reNq5hnLy+qZOOnSDSYX3bYQi0SV+vADG0Og42t7ue7ec6hLSWoUgqym2P+
VjtORLQyms2RxKpdYM/1EdWOYu7ZVb/hX9v+VMvNfywMh2JuhFXjGHfZopRU1NqBFb5Haq0xBWsK
4VQM36on+HYzF7dcxWCqyG7AJJTl+apfwUYeBh9v6r985M+jLDK01HXQvkGR5l3nEanTXPO/F4/L
D9iMiG8EkX7nsNJ67piz+Y4mxde9awkUCKpJol1MuVfOXQ9O/wTJhyBoS9BrPfpKWs+kQVkMAX4f
JzmjzYUgN3HnQ/pfSb3/B8pySwvubyvrTUfY1w9zW6zNDl9q/GhGscsWnQNQ8/hdaWdrF8E8Irt8
LtRwuZ+V5O6RUOvKC8bxz7CJn46rgUcgmDtN9tsyRifVHKg8efAt12tNyB9es/H1QbkyaOPFGag7
Z/U44FXB8e/QuimarpoAj6Gmdo1Q93sBjkBM8WtmT5hQyl5a5qoI46YisXjKOVoHhJktvh4Xu45A
H1E4a1DfKbLQH4uMo34is/dBpj2UX9ehqusK0/raG78OSppO2IZXYWuxDOCtCnvtra4/SJ3mrEBN
tlIyH4rJUph77/0IQdRV/pGRr8+Evg0FS9ceSofRxsaYXtxaEJaDr0wzX8yWsLAlVBQKorgBFLFR
2uWidsC21rBw7Je29iThEP1zt9zcwfWFnlzcEUWA8V38R62siO3JREjHoOSPMgczjgrQsUgAFdD7
9Jss6m8GAGgzH165c27FT292a3nPPVylGcSeIXicpsvXqbeOUYKY8g7s9a3KhgsaqX4JA5XsFeQO
8C5YEx2rKlb+llj+wgFrQ4YH9gGY3HgwU6Mo9/gxiqViFxpZ4Ni7FeI12qZKEII9ATfRDbKpArGG
6FF8bXALcJZvAMcclBWMfyXbkPysL9XyL+TshugUyhARNVldeg/YMSi33UeP+OQmoVya0Bze4FE+
x42ocYpyohFWEhtf0U7laKRgRDl1lbcnXrEG7ikyuxMR3FjWLFSj2SWLyOFSRH/mclRGD3FTIn4G
BgkFV2DeJGWwjXLJ5PQf46m5E989idWiVRtLpKkeg5WL5PuOwB5LM/vVmeAaRCbJ7gEc5UKhaZ0K
0YPGxt7/k7qfg4u2t9gDNhFlq/aWszdGCZMd13CCgHLs+XBJ3tfKtNtficIGNVdbIS4Ezf7Iq/fw
sksAnHg8dBbAxQyqSRq5k2zb1MykHuEYCGGkIrbEhYP5qN+fj42x4uiCIM2MxSLbsbw1cuhtwiVw
1EK4OWu/lIH6wCP6yuUG7+vepcMaj0hxF0ee+jubH7eMAdS546dQBHZ8MFgF2YcLuE1ymS7HEY1I
wAd9+PAn/as7ZW2BCt+bWc4Nl3d9Q9nvEt4W2n5pL15soBAvHFha+lh50Gnra41el3qVF/6pH8FL
VMqypxjJEU6awoQjutJheGAqhwUZHNC00zDuNI+v7jTHHc+J2N7BHbNJXIftgGSjzGAlB4iPVf/b
zmaI9mIK4ucUWz/OTkPbMV4xVMmt96rYbF4O05MPAenbGhRVval9JFSmc35ClQWmPYfjyOnohW4H
kQvNmBYPh9QGUj4Pho8nyhV+M+MKKAtqHIPIt5X+cW59YOifrW2hpqVzjhNP0kQdUE+OsOIj7xcx
mJ1FYnDfbHSdE8Ve0ae7Riyz60f1oT7zGqjSNgkIKHtSBKzBXAUrxdHMcIkf8/muVEaph+84fjdx
mPp56hGIqSCt7W84odbex12sPErHa2SllJ7TYzeO5H9JsjXd2CSGOyqAf9tl9JR9Ay6old2Xwh5g
Sw/iOe0QwlSEsUdtycLCxT3HuSAibHX+lfPjGwu4zOLiMsu2SuCfKne+bk0eP5oikgeCpmvAXFRP
TeiTJoi6FFoj5vnx5MrFbEMQ21UD/yNaz87nu8+s8ermItTJdZfyC7tFy4Vz4GAviqXMTzZp9mHd
PpGGOCLVmmvSs4MZqIEcuGC+uc3M48hxq8pWC5uJFNEbmGjnl1pyNavCOIXOw7thlVBzTqCUMTHG
LOAuyS1JQd/4d6KqSYiU+QHgUuhrHeaRb4KvVVdczeeD+vudGdHUwL3u1+xCTBYXjQJq3f6YnfCI
AC7HfZV22HgXwqUo+agpG38bILaGP1Lugy9nVK/97YMJ0BgAXH3V6swrhBB5Ow64KxmALBXEsg4c
2tPovzDf6qOcq1GJouAfTUlXgQUW9QnlSZZbOtyxYW1l74UFUKsMPa0KlAxOh6l4dIO7xxoy8RVy
ZR4pVqlngQe8EOC3WDCQ0Nid+NqJbWSWaW1uktDMzBQuG8f7ly6kfTp1sBsABzl5SOGPLZcNwCyO
9R8uihME0iSoatqGKYZGZ9zwsFaUmK57bk3ZQ/Wlab4TFmLEjKaxRKQjSOSh3a8f+ELBRtrLbp8J
OsHjWOqR0DIA7Dzysi2pPhPXGMl2wR56JMujkuTtfxEhDPck2U0m7sJpUMOQsow3KS/RaoD65OA9
ZGzrPsdEI6km9at8Zt78yzsi5b91bST1G2cKnSbSwZU4fq+OFIKJ9wkNctZZQ/DXBMfaveI0PJ2M
LJiBHcCuhb2Aefz9Vo3jOJs02akV4oKG0iy49u5gLtIawZCjvvK4C+Nfzy8Fu7tfG9tGqc7Y5YGa
4GXkFV+LjS8QTpTTuB9ql8ZOH7fl99mHikdDwGWXWWNTMY11uWUY0j9TCtVLLn2u71TSMCLHLC39
+Jln9e2fo9UJVAJQWayg8mK2ddrmaqoOUT5ExJzmC4TV2t1edTTkAnAydgc0s8Q4ppv4lczKERT4
VBQC5LPSKFnndjdArcLyPeo/3C8Njotf0boQTSSHohzUT7uIAigG6aAX2WtM4Q/bAKVOPNNsCMqa
fEnFnNnHzEmaYxdsjhxpQWu1ynx1sY9mqzg8F4ocw0rdafhhyuWfjv84olHK3M5s2HK4zUGb61Yj
QTTNZ2SZ1XXY9f8DtiE7cmhAU0mWNIsPFJ805ymj/Q0Mue8il8LRgvBDQ0Y2wwll/G6GQ1WLdHE+
mZIcuDXnSjr7o+TKv+atjJWWqoRd8vQnVrnX38aoSvoRMLrSnWVXigllFN9R2+VKyu6NcT0C3EfD
s1JWjyltkPVnBnKb/Tdj6NRQKs9DwHN1nTRRd2vQOmniSnpbnJDcwadVF/7UHnxK+kZaQkooyo/y
d7ujKitZDs8qMQBNyYvA1xo04Y0N+rnJrNC7TKiIBx0ulyp6BeRSbFgZx4fMokB2JOtA+DKJVtVP
J4fsqA4mqTH+u7N5dsaM8hMp5OyJChYdneWXh4PcxJh312CrKT/sHUO/lUXuF/mv2vgWtUVTv3VS
2EZXnQnjnFN/8FZGNuAOGHUivXnRXpnOcbBC9WQI+DxatSnAYPmIDdJi/LGgR0RhZW1c3ineQ4O5
ve4xvETOFa57bjt6ap58poqltkUYkX9dt5OOJNy/mmryWkNTXuOeF4iqR31LotTerX7SmpOGje3k
Q45QG/7oW/YefL9NtBoTK34pecS6iZEav1MLu/BtAgcpFYZfgrBaEaVOan9ForhPn0FUY+2Boli1
/4DruLQutA420M20WAMIwHBnwTsoMizBd0KChkwuR8cYMBNPgKHuauS4KfZ99AY9nwF03enWaG9b
iandxblxFsv48aeQx8Yj1PVTrkwZhdz9QvN7sPATxD+XdiNFnTWfU43a+TZ37uHrcMkqe1azEhiB
gwRQAfJIInwPWcZ7MSS1L2Ahhk6X6HVW2Gb88SNFrhOpU6lY/saPq4Iy7U6Gr2zsFf4aJ6TRAMuu
Ma7jeCPNsI00TXruKd5sFwzRce+Hf0j09iXdIm/UvZN9x4ij1yOwgxV4Xv0iVZ40uHCVTO3S1Yeu
xuHTAVguyPXukcwk/Rusuvod3dr7v06pIHKjgHf/U/0ubhUkMT+CFWtt1wVuSXUGDLT6sFZ1430P
QLGPc/Xo3iVUG9BfQzfNAn9eizxv1whOx5DSepAWDCiM4X0+herhLtOAVq1MYpV7+XZBteBq7V04
h72CPI14124YOhuoNh7lNQ4LUS+PUIQEN1fXkTJrCZ8vN8/xdzOf29MRHzGcXcLTMyu/6kC5/DQC
VzxrlOLAIbh4vqCGKP8FdkoVNB+oTe6zFLqniw9ynJoTnkWYkQjSR34iIbQ/FU6xzhSW95+VE7W8
rSDGlnto5FegqEnCyxdD5ANvE/hmaETKzC1C/yf0yCeG8z9Qg8FaWUgVK3tYGqgksbWlO6dMBQxD
5NFEv6gFmbgIMr2UZiSG25YeGLtoK7KZ4rVBwcFdFykNx5aDWyOl07HaFq01CFELXgshVEPOEVad
tSqTjMnSPhfKLILfNt5zIb88AFSNlL2tFpF2YcF8rLx9zgoZ7W/Pk3Ke1mup/umeu+zLT2ApnMHX
ABLRpX4cTyZj1M8qCWSLOBJWaLhgaVTbQ6tAQANBHcSEb4gzIuJhFwD9/QoOxXvRdNYCGV68Jkik
gtYni74VHA5DQuh649yzSkAKWByfWKev7/r6/9v+3ZWDUDlB3E+tJvGx5AUbzuokC1URmC19DVbY
H/fy283ZzYECV6AQvZ5f4yJ09oqRUpnDHkEPJeNnW0lnBH0lrsK2cHEMOq1nEWgZ5OHqFsiOjhnM
BnUjREL2dsjUw4nI8+Scuk5bKhjsKhJEtspoJ1qbR7MrPjYOnvYAR+/buiw3ooy7gbIpE/ezVE1b
gjii7olkVvVffqUUJGnZhQfaufaRoUubUxnO6jFOJa+mudCGELU/r2AnZZYnHyWnzsquAxac+l6o
61ZSeC1oN6dGaNyue5a5pGCBbNaP2pjxYmXmKnqRJcj9LrBtKpVhQ1AOvsma+YMhX9KCZCNmGbaZ
TZ0U0ShcUlGsNtsrKrODYtoqIV8krTWEMFJnWrXwQizs7PFV2d9U+kinqVZuzaI5Fh/x4J8Y9Asy
WT/8p9iBMeaaOwD1acLl5RqLjMcatdcW8uoABgHPhkezm7SwxHI46TsVulLjrAliUHgbqqXKwqgD
jIn6WdyXfywa/H5t16v4vj+Lfwk1LgGNHTVvW12imKMIOD/tFRgqS7dWkofwRK66kXmtc1BtDNep
o6jmUixn/dhiafDWdNmGQJqP1SNb9DErO0yzdETiUa7fflvzfyJ+Ki3t60mT+10rIeDHSOoa+Fmq
n+SA5XGTiwdQLHv2yOohzW/X6/asm/J/HW9ralzgGUV2gkT7IKOw+StwjfWxFe1XxfEVPqUCPv+Z
/6NcZT3P9AVH7AwOE4JQ5/3JokzhFX3WD5CP95wjzXnrIGzqJ2Nhl+zy8jQOGM0G6GmLGlRY7lkX
XPcj/TV7k2F1DFCzX07DWyDyGC/+xD3jlHkDlDSl6OeGocsVwabwlI4AfMw2lD6oCrLhCXID3GX4
AREBQIajbkPbqBDLkOLUzbzTz75ZFseiAtyt9LvynzJucr6k6fDXQo7EMR69nucWs4x/HTpMF2G3
RTtdVzun8r0KS/qNYi6STEaWCqcN5qLHngWr+D/CmbVg2z/IWBeOjGIy+usmpI4YoyKwqdEztgOc
8OAHT8tW/u66j+GWUeMR1WIgYZ5vbw++orjeWA8RJU2LdhnsYFQaCNrhRYj9KzYdFlktA5ulDqpl
k3ZKctWyd9GqOkzUbGaujLCwg7s3LSxhmeyzO8zKL2MIPjJzHNr6jZBUU6QBmIt7muwKHViOWEVt
PmzwUj67OvaI6DHbjlibPqMzzSnBqkVh0ivnRBSU7cnerZZvrPc7loEaTyVMq7181/hHjhaTU5mJ
ZkTRVxm7M7EdlJq87LRmPHhR59iuUI+WzE79xfgi++PovLGHSccA6OzOXN2SWvEo33OWNixxNWMc
Vhs2youh1lQHI8NPLlbAmicz7YpfGblspNlyj6mk80nrqBkx/MESbvtNA52ylfeja8UNik+hPSyy
BxWFBwS6BinV+NeTevCBafhjNjsLJtTXUc1vp+7WIFMtXiVJreQReVHQmrcm49t3j/KZWs7Dvseg
A/8E+Q4ya1jt2niT5+yOhJO5nj9LfyZnCzsByLzdumffEs9VVzCsByY9aPqr0ElBQVFEw5Kqn+mC
ghA5hkzP1t9I5mznRjI8OdZtlbK6sxtAzZLC+tt4NVjEA8ZS7rHBh9S0LLYFIyD0bqEMMQRLUWqV
mFHrrb+UBA14F3AgGP36+eBimUnSX2ViCwvUVviID0ZCzA7P18QqwHlFzo6zlNtLV085RlceXHk3
0zZgiccIHv+GNy9AvZiLMY97R6KAur2VDfxuLkKdYLX3MjYJR8gUzVshlnURek8ECLA2wv3YLU1s
Zxuu1DJ5xId793LGF2Khn70C3/uEYXp38ijdGkQmQS+/GL1zOpsdxLyxRxUoE6OPK9ub3+yWHJ9f
PLi4CvdmjuW4b7GUTYj4xT6SjHy7fspSObS7kzyNoHDaVyG9vnzCzfesYSr5h2cEhy5BF2QT+68M
HFW7mSyu12jhsm+yH3NrFbKD0fmp2h/4DKFK84vq/Y611KLzxxplelNEu8J9QLJdHn5W+EzS3rr9
Jb663YL0taa112Q0GQgFOuivDW2nSfftRLMnR2d3Yy294DOWW5oLa9K09HLKaHToeYO7aL+cQlo5
SyVbenUR5D0TvoVE1A9niRm9uWY7HsH6YQr0x/YLJ/AoOi9SDbKuDwNzq7Kd8isRdJEQQ9NqCXxS
oDydGhIDZ2eVXEIYhJ4ySkmB3DV31v7qTRyYQLAyFnhnh6FnNbHv9qPH8G1PofyR5WWETlNjnduK
h+plbx1qtpd88havCHZi8xN1yyCuyhYnZTHf7WInv+W6yH/xzAcXmNgVZpPPcWgMe2RjsMfUcUq0
ISBI4MzkebmyuU5Q2CKVRkTx7WcZeFNWrOsvmXrS0hgsWihn1OkBR9D2qZ0Un5De1lfRR8yYzwcu
M+4yy8ky4k4SgkbTYOSwcbUE4yiOTMkgeJOqBipRGL902WFdB7dChy8MF75GCj1YY5goq9JaBvwS
ntHv0cbIz7RBtmva1hsYc6Wto52LqJD1z4i9xDTgNngfLBDyBIl/e68PRtJQTRTt1+AL5UE/6bxA
MQvXiBdvgw0POV8AcGZ0+QlJisQazGvAx1R0CA6pSOJvJWFF4dHtwASMGmVLrM6SN4LFt2ZDzdNu
jEf/g32wgIFDbBHBbJzz3/fl1rXSuA0R+JS138pkK7JS/meaBkVC/40uuk7NafR4vy9qLNizXcyk
ncWdcB3pDKBheTE1NVVdxMLtDIS4iYDkdfXuFDQw/uO30SxwNxxfumVJFvLeV1OV9KeEJUE7MuYf
uCzBn/IZCubexosxncrAWpniaXxmMazG6tlxbbJs1vrv5S1MKWA1M8zle/QWN55H0xvxvKc1JYbU
nQ54ArWimWFloLoW+VWSOx9GOIvspewcnJbNCLOjkRD0viajjsdpkBP/eGvQHtr+izYiDZdhShW9
1TMcz+aJMRUUkSR97DmP5Ffrb3TliL5Ya7hePePyEaYFJdo/cz5X5JEJQAX87ioQzs1pOR2IFWIC
3oZSezroUm3SOKm9v89qTM6riIG1SGzaA7Elf3oJmldH+nQjlatkEHRNDw0NxJwOAAo1GOlIiols
ifGlIKuDkZHGzyJT0t1HBSfWM2Qbgb533t1vFX61fPB+qRRSSDOxvN9Iw/oRXhT+78/gb53yUB7B
0WBuXQPW+w0RbQs3NU87LSkALoIA2rTgAeXmOfgDhrZwdyDJJoDbIF4D/weg0b6nlTVr4+Ig5/5z
lT3ToSfP+8wpRG9i8r+YUptU7ZAJ01WGxYs5fXCqryQeP1v2yVvDjqoRSy0TX8QG6Zcn5sNUsJoY
YVnS7SUK+LNRuIu3zPRRRX3FfbxrEZdCF8cmLaxxJsrdy2rG0jkBXp+TBUSh08buL9dWgl7tYkX0
phlTbjminyadChpo6irKEyjyBNBNJ/vU6dxv2e2Err2tGZEFresOjFsNeymL1iYjSfO0omX2L/kX
qvJptg5oDiLOjPKgxYOpAuTDpiCYU1WoHaxQhhy6HDg4TMdjZe0VBkOdCRMaoyVJAnvCg6s+zvWv
WaaRWVhJ1sKZuIJ+IK9KyFM8pXHdtcE0gdbXtIJfhUsuRtCYa9f8vlUeOsBQFDrTtbe/Cawl27dw
n8gNFG4RdjTj3wFgooe2RRLu4F9DWfbHZAw/gpFQWrJlf80TqtZljb2okn+damp1Z58eEjgUOib+
w5BYz4Zy7L7TLs4SdWTrpjonRHY5VYEvW328sP0d8tsgn98cUlBcs1TtnyBZbXOqJVitq6+r/DXg
oh6ng3FKfuR+jnzM5uxqdoP/UdlMEtaXlrISOX7hISv6F/1Sjn/9eURTdp0EGWFHkJRCnqBLEvW6
PsIrrhefzuO+U/UjV9qbtsLQuwoiAuEgtYjX4jIn6m69QwyF1gqQWZ5ZeBwRdkLN0rudbeKQwKhx
6zjue2aAeVwIi5745ERi45ecWFQN5RU45l61KIkSpOL8D9L6S8D8xQoZqLtkRTO9xF2zVIDCo6hx
yAnLoG25V9m7xc2EcFVfMIWImhEdISr015PJa7XdS3erzFIc3PLD0bt36ohIWzBViUxcS/acbYNt
O3tKpsRhY/10NIij172ZtjWEgGeD0F8sCXS4/MMRqOpjFToMfgiqhPD46wh82dvjM/JjBPXcFoA7
Zz0p9boJTalVXmUvE79EYDfh19ozz+HkDwpn4sI9URcXGXwD95cvPTK/rnIY7TwmHHD6eWlVn4ht
VOLqsa3jOLtGCg8vS5oPhQ+r0YvbfYytM61+mF4V/f8GN0dZWktOfPyKZqceOtwR2og6h7Cm22nV
5Ux0Q4eNSFdTVsn8s3mPDhWXEN0aslrwqZ6GnHsaBULaBqen1Whm+HblU285CARreVZ5tR9meqlL
HCzWkNMhQnJDzKerpiGXnhY7BlbVkuQ/rPwTA7MEFjcmxi6TI959npA/I0g35GrWJ7CBRzasKp+k
8iF5+aKta6SnqZWzpOazmRKHefkzFlY9G6BqaRHZIzI951aY7h/3+GKMEir7PWk/VXD97PIOE+A8
AVMpbXtfCzKuni+OHFKSNYp/6wa/KMmdeDSWNUSON6yq9AlcV7dyQOehuizxuLPxOWldRw+8xDEh
8QFtdmvKi9PrvrbSoqPzadubCGwGUtQ3+aLGQXwhS2LYatHwZ0ktTVuYhc4FekUGaldOsmGsNYxh
5Y+EJyYwmEwz9wLSXcq/HsVWk4oRI+aJ1a6FiXaq8/PbnmuR8woIaP3CGUSh/+YKmfWro0MCKEdt
45bG3NpfVjVZKxJCnnS74rZZMmauuNRIhRacFAiB7rirHWoklNQxJXc520D7JlKFZc0bnsNwpDug
Mvu5/L/4XsB6Vwn9CaeP45CxmfFlRD2YD0GriK0uS/7wdYVd17fv87Zs7AKCZfRvjT4MjongisnH
GbVyKvIXFb7C4B7wjpLsR4B/i8IoTeCqJImBEzJCZn+4O0CnsWVG3dzM9I+CpwXign2CVXtB5zSQ
WaW9NFrkqFsOnlsZLlF6UCjw4I/xw3gTNHPFENV0yYTDeo3evB2qXqvQbQgZQfn2OId1II+IpqBb
T4d5uBfmc2eAQAgVdLNGIKybS68BfVYwVlH2Fn4o5KPcAuCVA731W1iEgr6XDdJo9b2qjTFP+viI
GyCptcgzY9XGKS6ZtuiXft7AphkAMWzY65bgr53iTQpzYfPxi4/GKzFVSSYGKUvwNzHQOR7Q20sG
UcXhNWImdOGaFzu57VKpAHJnKImXN8j+F+LJt05mU10yOJQQKuKZJuih2vWBMRz6BZo2s3T6v2Gb
Tm4ewr43PZLf04vrSm0xPtx3HZdxIyj9EadfiXU6vCbKCRstGdYNlYIfU1z7JZ+lY3MzDYiifk+q
SINp2GolLFwYnvBs7H0lCXPtiNf1vA6hSEmU0qo1yHLoizAQ+9a8aWM9NaZAc1U0MfqsD4FzIg7/
OwIoNOJ0b/EZMWVGGVIA2r6uqnQmsOD1HRZ7tzMPDEJTCXDG5OiXjKEHWqWbK8CliNX4b2nL68UF
N87kkLqqsEIbHD44RvUod3eYGq1CgVriOJCeTcXxYY6z2/qEGWmcp18ufExzo4jJluRn3nCXi/hQ
AF8zRQ+LRWcraUk7Hl8qCl+A5KT+xyPhnv2wNDz9HQQ95Vzr+vv8PNV+Wp5s7ypm9Tl5KNDty2IV
wnDYMXlguiWJpBVpbf1sCdGDejpvgW/AbbEzSpXIE3lAg6gGdv0c/2vNRHEd0BcNPnKN7GjlS/4/
N5HWlhavS/FFQ6OV6XuxuFzh49fwedLIGrJhmsoIJKv5dsMiaQ9k1uP+47UFuYTZDkUTtFuVQGrm
4cv/rzzqV8urAQV1uMlNJTN/RPEO3nDJ3gHXjOI12T1/FOMjRfwF6oT8Ppy351iIZJ0WkoC1Xvfd
2LYrjyOklPVURG31PfyLxPyh5etgOZ1RT4k9LtO+nLzOzEYFz01QMXiNStwzoqIf2yEdCsupTFG+
BsFc7HSTyTGjEFpU+euUlxJYWpXP14zQiRBi5K+XfHmqXRPeHWFlMZf9jMh6WWH/ZJplDAKV3NUQ
dMdYLeTW/mn3RL8s8WrlcFhDDv3T4RlsNMlNlDoUypE4MiomupOnubns8vFbS0L/omW8MPBNWFZt
qY94l9xWo/FFihLEd4lTkvMRd0Vp9M6EADdEbuUj6HuYcZdKZQTv82IDLdWofcogwAZPnNLRFQAK
XYYPb0gHRLGvDQHc8Crvqz6MBsJVI4YjlyKX5t8a8BUb70TitLgGWgSgl0PKw2FbOS2lLpuPjodh
CxVvLDHjksjxWE49qGhUQBmM5mqIjfsKO6NWTpKUs1CyZ9Dq4JxQ5tk6+MdmVvdyBBGHimrS6x6y
RWetN+EQwdsOHIHjU0kcHN2KjNBtEi9J4vx2ppffwFDaGWogxS19Ncg7rq+k3wBLhEdP7nK4Gnkr
NBjWdmTOm2GkUlTOAe1tkywUVk326KI3XyujbvZzNjGBOZaMBQO7VI4oBPDjkdayk32FZxruBSDZ
iYuUkulCc07eIyTA8MMKulwSW5f52kKzKyr6H0wg4N5WU7N1eTnog4rzWg+neZMhaB45VmRjobvj
i7ShVA4oEs2uuigigyDGYODjRLnGDgbNlvZlfwUPAkWcKkxfXlMczBwUss3zu/1QQG5jTke37SYP
BKrb9nDVUQTodZmdkXb/UaJKY7/mFVUfSxSAG9FwoMNnfEbwlRBaaMGpobZwRk0EB8GlAI5jjn2h
BfFC9kcreYkFpOZhJcs/BMcx8smSijUFzyDknVMcsj8IyfaappYYE/GeX/a5OPDhCZHwqNYKcjqf
kTVF/NRGotzISy4txuS5b70Xd2Uczgjqg5Xp+r+wbSQxXd2zhFlbsrQl54jS9u8vFeyfC5HGUJoc
+HodCVTRd2Xe6eY/GYb2s91KyqTAi89a2/diY5cTZAPijkVXHV+AchmOZd6KJI5ngR0gQAGKw+LX
QlvfXFXnasISzilFY+u5bqMrOtIgvcFhEkAjeYc2nUFS9EvCwQ4dSffUddtqJWIDXtt8DE4+bRt1
y4pOdrcia9+MGVn8ETd/V4CQhd0rn8rHQmYsQO7nmN31jk3kSidLi6Eg5sWS3rOrDz2WYWgInBP/
xsfOvQf2CB1SprIbE8opRF8g6y5YJYC4RmvXvKIJhLBf9+QzuVjoZPxoEYTpyyNvrGlVZrLJAe5z
W4EVCSpv/lQCE/oFYuj2DMa7Mkc+kB49toiHAEYehFT/rPPQPY2R7OvwH40LMd2quRlrRX/fGomy
sMcA+Mzdv084XVrSROrecGSidW328xrqrRll0M9xgy09Ws2wT0wq3NFE9Y2IYnp3zfysCf3onN9u
Wxph3lUsfoLjnwyUqw5sCdy3KUTR0KYHqGOopIQ+JEvsXOWjvFz3OPS8V2PmckBs1LAppjsjtfK9
dfxSVl3gY+jS3+jJKmT2YrvxNP2iwxZf2JMJ2zIzWAGAGiK3wrlH37eZShY/A9r+ARXf4TxL54Q5
fWh+8NOdWPEP30MdMG/7eigAUqXDhk7Oqv9mwKSsirxPufT/3L26IorpA9XRw+awFHBPZdMyDRMY
t9c/eBA1bDzdYCUdk1wp3ca+L2Tjb58+Du4kGm4ixFU/aBj3yKM/acyXJ7RJerWD2zCXXR2pHctN
p1K5fPpf0jWIGgI2RWaFPCGknIyD1J/aWhO06sHvRKkxDS+eDeg5bIrxi6FCRgc7wL7mE17p3xAi
pvy1c9ZmmL+/37gY66fogwfjudAQG7dtF1ILGinOeu2BPohfHRfHcElRvvwpXtiLEyqSLBabjw3X
bd59yA3kgwsBcGxKfofJLMjFi1Fai/5JiagJGAxrGBhtqEHYn0z5XjW75PqNeshhPqxUwRUFSElJ
hnd+LHqvgjSljvD/c46tlMntX+WrjzR3DjJz8cRFSkhHN7I585mbFPf9UExgW8AwCqnRJIuBec68
c++K7J1zQVmNqa/jwg/O+8twB+EeSqzv25LdzIoUOK+UjgmbntQt7BcJPFLSjVLuBQZEsaYkBoJb
u8nBsmVYvMU1Fg2auodjiYtOEBD/VLJ75tHtm6ws5sNxfavokH6BVQERl7pNs+6xc/p9ligsjlLQ
F0+VBZJRUZAEB3HVYybtRDsBpIcEYzOYbzM/lyZVfK8QmCqDvMnWs0FAlDMIpCZbVhMe0NCfXNUU
0xPZS0VJjBc27Q2s33yupK5eTAawJd5Q8E+OOka285PbX1+ik0b1c7hWFrING5CPalmI77MCCmRd
M8ph5Wj/8hIsg2/4Lea9d52JAmkMseGNtOdhXxNZZHgWU5K83AlhSnnnlULVwTKBQ/SzJGp3pJGR
fGBPSLlL5ePaUo28iMKb3WDNPRG37cZr6DmeqXcw+pRsVeW7Oh7A8nQVJ8Vs2jRArkaRo4lCPqBz
6b88cRImToLAvJEBy/uLIsvJE0QxzYw1DoegpWC609cAhXUZqRb+2PdSBHLbCP3igoq0Sw1WIJF4
odipWnOXFm8A42Jd0kjI4YLI1VVy+al+pZT2H3osO8dq+PYOeshkDl+uZA5g4SIlSoclED+ihV2h
JfI8w2xwiGKsP1oTIdk042RuKoeSCR8psMoJzJ/D6Khzc0iThR9U4W7a4XQn34YkmwsMy15wqe0C
BRt94qzfHqeJwO/6dX/Q39WISaS27emGFnXyDSDmsmgM2Rhi1nzMi/xxkGQD5MyrtiPmDBoIqToB
BFcsrkyuRKCv7Knhd/SBI8fqonRzb9R5jy7QtPlp5xOyMM2sxrSIAUgPtELTSAMxB0xDohYY0dCk
uz8AeGgVGpCA5S86NM8oFl17+lBHS8AQkoEGneyNuwtgY/N3zDOym5ZDtnvPVfpqyW/b+5JB0X/P
U3R+plyUpKLWHRL/yGB1uR+8/GIrz5SRHof8mvIwbPn2OukgTlkaPaFemtB5ENXA7B8yYMkwTRU7
U2Lw9f5wo/t6MsYS1F2vRMQU4si/FjKqZ9RD2xlOq7jrbwJwQFdPBpNP3Wi4BMzkE40F8QNxJTfX
ExVZ1AR0eOdFjF+NF2w0y2CEx4OTOIMQw7BcQqMIS8z3Hnb1rkJ6U3wiC9eLMqJ7ukcKD4x3wPGa
8IqwJawFN6X601qUSOTa6HBj9iaD7ppUukJn0DPIJU1PAuM7XrwgjP/ZZly8RrcJwCvjxTOVKqC7
rvu+pyqgoKsceKLxcoqJe1tMOeDoQrCJHmSc/lEF56KA7rxJQMtQ3WAQuLc3RGJSvEsXMtXi9F6F
vZ/YKqGMwT40+XOWUonFsInTzt40+fABtcD1XJC9fS62PptmK4kDAbjsf++zujItXRW8lz08gEc5
ZXJ3c8SdW/5sEAm/1dY2mMePohcz5/xgfgYQjrjP0woIxLJD7XU0ZJnyRGPGGaznmupb3pXYZe5O
ygb+hqCBmsD+EEBZJknoauxUQtvGljUoTGVq+epSC02ynB4AXS26bMf531KfdglZDbOQTmQ31mto
6PTV60UxOldLPe0KqU4iU2mWW6VBnB/TfSES66Ft/PWYsKojFCqBzIjEBvGytz3CLShetBN5Z8NH
+bVNyuqF6J5Tg0N1BtpGOq2E9LlAlsBDiDnxVZW77LMVEmWROU2ULIfGux/D4v0E/yrdsmygOQG+
QvPpRMd9akU5AlsnCwlrVZNUqkLIKowzGsaPeymlsQ7hZTyeM7Yjm6bMKLmEJoTUYoPEZ1jTgxvh
YLD16t7AJ3Vl2ZqA/zxZdGIAhWR66esBBCsOYHzRPJ916aRecFM455orgL8Y6Yvle/OmJNUJmBDC
2i15U6Amm+me9v6mRxZFp0qgSnDBBnGSSoU4aYBWN4orTTPkN6d5P1V+fgfG8AoQABeumJvxgvZV
WUS9ep0sYkYZT4ulUIxtrlvwZfstbNuBEU6hmpuH6fMEdREmf8Udu2gPkoPvwBTWkWMLuqf4jFs1
zFEpgphC8NuaZtHFfYOks8/IAD+0aEI9RvMAb23VLN0U8bN2+ZWC9pC3XF+CDoAlz8VuceJnDbY8
BxacmXgFiyJCM77JMnLKBeqLsNtzxL6xAqNkaUT1gzSB5+R6cRb7NJ+TFZ8gy6ZIREQ+0rkDueU+
Ls3SDbflRI39crstd1mPPUYmEgYALqwXYPz3pOA3GsAqT4WIQNEzSSlsRVUpOrmKU87aQeKxIRik
PlWGWXgm2dPQZ6mgFW79gFt5QCFrl/1mRkvQx8BqCCdeydAjyJnGjz66uYRbN0A5UrmJH439bhTz
QUv02oxzQkDOvNhnbIIMAU6oe0BY/7TR/Sl3Q8GxMPoFooN+uBdLwq2uFiFWhFdVIQIj/FivJs2O
t2gZ5Hkyu/PPOXWiFszxG6zXIQ0nsIlgOXxbk3NyhwAEDwHU5Wad/kXQt7eXYyTIfvUJH1uT4MIk
W8UsVuxSDuqZAkXQVCSAFevm1wovc9ZMax1B4Na4b4nbr/a0aA4jmhag9O6Z3cvasKQnEm+pw7J7
QtXlejdv6/XxNGIUqtDbiC3CTZD9jL4u6GFgHLPYFnSYYzHFFEqSx6hiGgtP2xGfQS/Nh3jOKKSE
HFKPa7Aa3ANEjyGuvblBKnpq0/HgEw4REGxRaEE2gqrqw2t2gvCVO9ktTTm/29tYu6vGKpAkmhu/
rf7pYHfYT9xsACVHpB61TeOLkAWo5nnnfyYkW3KXMnBT7qkbSKYQ7mu1IhvwAnX02bJdtJcTR/0B
AJC5uKfxsROB3I4FifjyOfmL1t66wGxeVm6Qgp7ydE0ZAInZ8ykb4PEmblDaTZaoQ9GEpt7UnS7T
aDW4pPe1oy+Geepsi8whpMo5Kury3ysHh2HoakriYQ0cgKuEZYbGE1c3uo2RRqPZ0ELXdcwKcx9O
O8yuICveWgGzTcS6QBYjRdAMGRgE/i9JrfE/Vcxupx+1r7Y0GrLVlMZtUDPIN8kRPBEZzbyrkdpO
RA27PtzoGEgSU8dE3SMIHVMAhBtpPJ0r1rROY2smMeoAhHMWGr19OIXakUK9B8zZC553Sc0pqEvR
Of5fRJjOknnbKJhdprpGR1Zb2ELx/XbdY93IXMWYkdigZVskStRf8zMk09xCQaiOYnfKpy8X6x5y
jYJGC9MRaCsaeWnTFL/2t22zy9ZzKlg2iVsyxWTu/xFvUTWXHHCKlCvpIpfqn1uRPq0j6mjexcwd
SI55SYkGz6QChoCow0x0/vvmpJNN6jI1Ou1yl7BuQMUmhHp6HMZ14cNQDwKqGN+ZgWqIxXs+Wbhg
K8NDCWZe0ucL+MnP3elNwMVhSojmisxGaho7lqHIHUD8bMXeTeTrcyjN4grMHDZhUQ423wpCefhD
yVhAVRDSoa5bAGOnFXNVTuCAUnaWCJQfaZ52OjlBmpZVNk9ka/uaKdrCJIyNsjSo4sU4AlrWAxKf
vrers9xfUA88BiJvcui8DOvB6kwoyvnuTef471bjdwfXcElDia16yAzelX1b5c4XliIq6dpVRBXX
Auas53gvTy8XRO+iFXj8fk+f2BUSvEoY8U0MUZ0QuNbdVteiO5rWMZSwsvpBIl3rA1AiWtXsSvdm
T/34EpInE4NGJ2XU3FzDIvd2YkewuumuNdAaKXlaCdlwYHDsp1Z0B5yQ4gfZsULHulEQXun1UGov
5kWGOaznylw6bwbxOaW/pgpTodgqbRKNU+S9zmZ2mIpxC6Z7ablmeX08LJ4JuZ1t4LxzAF1S9q1G
4vtAL+5kvS39c9cfyRWVtpYNw0djbHoWTshRZhTYWXHOp8X2qvaymNyK0c661Boab7A9IoRp6WWz
iMmdTmIL/DqsNJxb3V4RVKJpxqJe8s6kaNuNh6abqH+1wV78amA8jJvIbUJiru82x94elIl8y+1q
4VefKC/9LkyjR2r+KAk9USDDEHa1kB0IvbnkwE5EIAEMWGkcDFLbK7cQyCV7q9H/dSuXvoUg9pEZ
Tu+qL5uhw6CjPlOI4F0xhCm0s5rIL/cTpAOPww8Ry3/RsebI/C3Ibbqc9mSvtdifxVRzLHl8Hrxp
pEyaCGhIlnnhqlQ97pZC+AerVb0z1IIJyIl+ke49JfCnHOL9Dsl7V764P2ahx0WfSaovgnidz67o
UxHMcaMqEfbmxh7N/QV3v1y0Utg1YBWrfXr/B7WuPG9xOKjCHnhU6U9eSSiKn5xhBDgXe9G10zS7
au0CWouCIryK9W6dA0TKK31c2fpCblnCmtgRZRBXtVRcLKb7/26FUVg/Hv7FWbknescif3BkaHwT
15MrBwNYZpapZYzKMCzkZeEg215xQB7jivsh19witX393c04PjrsJnVLWdUmtYPkQIP5QDRdQYSG
chL7OzSjHUTvCTuBe1rSPIilzoJkoYiEgaBqRHveWlrOXTOtujrs0F4vwck9mLZqflNlxWmRXLMw
qFzN4VefTrqtjLjS2Rlol8BV837eliM660560lY9g8cv0wyqF4aI7UszBkAfsIQhEa166yYfUU/S
hI2T8gelwOgBGR882ZCpGcfm884I7wgroKMfKdVbSMJ+gk1OVeWeBM6ttFfL3rTsHwmxUr0wvMGj
V6BqbMaRMS+4DIxC/XYOGcZGT7QyUr1UtD5IMIg/H+lRouhQq7Cp7TiCBGwfHJMgM//ku50pbvoU
dJF59pbuGSET4O1ObAkEzJF+NbCeqX3Pu3En7d66GX38YXj4T+kTOOgF0bbRyQ67zk3h6CFstgun
hg/cGJbikLLYtJMlpZ0RvpM+DgThFIe6mUXsIEh/7gqH3En4yfxZ4DxfiZkXUYIViX0Vu+V8KtSM
Qx3DZwao2vpgbqcdN5B2Ih45YS8Wox755cd8c/1DMKXGYTMLwCiNcr7VFtFX6rmpTgi90pKI9/qb
3wC9mA4xNTCFssCID5TDuw8TO20mbkXPjiM089AUkv3lEzSpeEEQZCZHllTxNuCTVGgTYHWKMAjm
i6H4Epg1jLYVW0AmAP1KR1qNvhEuMqGkQTiMlq6dR9pFtLrDnSb7mTvqyLv4kNnvIlQJno/b9a/1
XKz13AGhErHoEg0iyeLuF7ML7I7mUOc5zj7MLLaLOclp3+Ykwwqg58zbDcbOGnylK0Vpf7VnjLpk
lxBh7+a31GV0yoCHK10BBonMPQNgVVk0Iu3+dzhPXH3dwUJoNzjfqIxP5EpmwSrdlnletKD/TeRc
/TOyRHH++uauHbCYLrlX3v3vmF2EAe315SvmVmYZ4WyEvp8LhUIqNaV+8g/0e+kW2kPV8vlnI2fR
HVAFo43GsZ3eJfXOhDYhRFyfwu53GSg3gf3yWfDOYr4foL1ETx44wOV0apGfHme3vL87wKm/GBR/
KDVK+YE9ivCWl1b/0BCEu5rmKIqdvpnz6Hx15MEyT9lMypTrAIsWvbPpU7iCuWUlYl1Ozj6nxSMP
6CclETi93r0mMpNhbbelqBz1WIIcbeKAqDSlokqNz1Ta18y52RD6waMLoPw3ED5qfZoa+4z21waI
soGaQ0IiyLaXM0s6RILvnyqt+g+nXVJx3qPye9/0nQLY5IF5ijpNkwN9T3+wYpEJHASx+7cVZkD9
1H5AwvyIJZ41fmMk1nQWSqroN561QXl3Ddx7/G9bP6fsvS+ndtPEs0jkw108j3kSS8tPCrSFbdSp
0uU/pQ4Gmi7scnFPP1qUpgn7QJvUx3DP6A+okZurHpdhrNJFYqz9x2jzZGKoZlK/LotHWZGOrCMB
RY58gel1QoOI3Oqeht72rQ+NSlnKD3DhVpTfR8W3kMRJcNxY/+LK3jAfAc2yRzR3GuyPTSjAnfRh
QVitaytWdpGEFE2UkH9/fo6uaQKkNTE3daQfiSjyR/xTMP2TYEGOAgOchAeC69V4cDh94uHevogs
5p933Zrf9xeZmFabQNDCjKHDwKAtBqH0jAxLkvmczvVReA3qpwaVZb2fWH+sPIm4ZVdHBu8Shf+s
wJwQGhU0ZNFmGEUx/JQLXKH1KKE8QSDhCKMitiL8jPYCkGQONvHpiNI1KKVmAdOF2dqi0+gaIFpP
ls5VWox919m5J60lu2AhXGkmdUfKyvl64sge6JCbURwfr3i38Yi0ukDFCFSjF1v79NPIFpDAqLFw
03cb/A3GFaJazVVFPjuJLGL63Dj1pRkje51QfEnJKgsE72j2ZSV8YOLvG8U/UHIJjUBvygsjtQnN
wsBFnLkjz7g+LWvpQDvpQIIS1weaovZqwK7SMdxxtlfwgxm1vMjBJ7iCswVCRBrGb6mx9YrGBz+d
39/FCbvQ8y+OVL1ntQqbEcDAJEMmW6/kd6ZnyYkjHy6jwKoa1c8EJFf7A0CiKHP0ziMFcW2tX9S+
pZE2cUsLlAV6rBsuzLNJB920oL6RxMjeaPxCKC9SXCTMJOfbJPhR112+lXRfMxI5xBxBJRLSz36k
A2HbXm084iIG+8U5B9TD0VvEQ8DxoxheGzYDSPNFxpd0tkqgjldNSxj6jMk+Q0Z+HGnLOHR+B2FW
5/H2wJxeP8qwEsPApmHCwUkrUzd0Sq/I8Pm0GviSdRYxQS6L7Hrnvj+4kApRW4ISnzUMhnGDjJ/G
Fk4Nh+hmntQvI7uqaqFGb/lLIYMttdgpibHudpyMEdjcfI5cyDJ/dmQzF949eWQkxjIkuBzt9XNw
9S/ApLZuWJakYD38t2ekh++3spbOoBFYEyLysYPpEPceeO5kbFIvB4hmDMDtnxQsvulVe463GmRJ
P19gw5CnRhvHQBZq3djNekA6gyi/P4pnLH+0kRr9jQwvJ2Z7T9o7d9LDjw/z0ZcAsnbGM2C2d2jN
zW/jiGMZUVNcVQKd6XP86JLvXCatHcB5NtSsiNpY1zfSN4oN+/QGMa+OAyzr4Wayh0u18NiFHkPW
fNyavp+jIRL+qwkbd7YFiA9Vf8VocWVhWMQbucDFHluXjFf8YLsZDf+1H07nhzKHGi29Jq4eNT4E
3ufx46FqpK2R9Lm1VAFynan6Q37nnbL8zN71/X95l20lnv0Juht4ugmcdBsLKNMWUGobLzPCAsDq
EVxu+9MkJ2nfztyovZEVrNZA0yA5aBlsOUn9KAAfoON1sPuS2qji6jN98hUvGyaSSW8PBRTDRF+Y
uoiphLemIzmVgf1G6lJIA8NOqkSSWlNVIW0PAPlx6nw8MHVQB3S77mKW2CZMRutUf+ec6H8US5M7
NIWh1FdGqWJ4PBzpM0iXX71VMFEWiCDYrbBH1YxDyRlyYcHJd1I59Uy2KKWMPQp7KSJGjl7AozQR
hGLPIQXE52z13kawXPsm2eyjPEKetfjJpgNp7sggmQalF2+fJglbY0ZcE5xuk2w5/fs8HjMV4nxo
XzK4wFs2+VBOUvCjM/UFCLTLIRZWBNdQGouIeP/fB0C1XXKLyfLo6tnfAf8JcbPvE70XDeG4oB+j
fR+v/rgQIaAHIudM2msMnf1LdOOPTt46TqHkw5W7a3re/ucvWs1iUvqsbAu+z+XtuVIJGMtznEVV
L8CcBeew3C4PyEP/1Uk/it4TEI8x6dUZIYbyu8UWsCHe7+Grv2V3lM6HgyjFapx4Cf9vC5fvz5Pm
jyttZWzL0vcsOV7qc7m3PQ8vQnhiXlCu/N90xhETL7HUzRjki449jyTjSclnatT4LXQlbaLtDi/O
elV6ytvcHEX+P26vyvNJ6QD6NGyiTxTAiU+DOjYmnPHgNHZPk4iy7lF1zdfwQ5bzpZmBHrCJob1J
xCV4QLDlVOVhfBrP2KwHlIeOJilPeOtznZXrF5bx5WwW55nCyQQEdUzs9CIXBpfFG2BRv+vo5g9A
tb62M5RDf0Pgm74OcLo/IIz9OuGGGXyh6f/Bk0lbdPql+DlbyNU5vITjBKC59HuwKcW9ZreQcnQa
IbFiVbZ9wxyjrNnQeP3cnVp5YIKSjuBfJpd9i1a8s8mTpoF9Rm4K4O4xz5/1udKnwlZXoAjSAOpe
0OVtdtV3mdKgCYXl1eeELzZ9yWW4+lziok65IyiPDR1Grf5j9CdMqLs+193fQ9V8EB/m3VENW/6i
tmkSQWhqOlrXJGCcHTXx8oQz+Xn5MkYmQUyrI9WPGqa9lB57UvFiIc2di2nTvdDl1D6RNe+UR6bO
T11RD4dE2IItGkCLx2IXOhCM7Kuw5zWqoIuG6Vy8jpfy9nuacbU46QXJqv4nJATKffdI0CNR9CBv
hQne2Mf+KRnf9QUSDqnAsuNvVUQ0dGNkKjLiE9oGsu6819pUZiKhTYqVQL7SRpI8r6SFTLc6D3Ky
lJ2E/A8kT0+bB71j76f5r6kG4JgKGlRHby/Hq7Ot9HxlAmozYFbscDX8A+UPIa8iwv/om7bpo8uL
kttyLxThW2q8hJ+AwLkdjYSCdf/r0nlyIPoP0P3b+lnVuqbbWaJSaBfu9dJndqNpSOQyiJbU4eUL
A9RXCvNOk6kXmZMkKh2jwNDKmdR6hCCtAzDcLMvBsRS6C995592gh4BSid4x4DcKYdyRGmz1Vyuv
VVFafIDs0HSbL2wKYW8DbzAioaC6Kz8raziTglrw9GUhD/zIJCMvhiE7y6fkM3mXAFpqP0Mie4ft
yluIHfyQFd2sHV8IdYBPkb4BVsmOfiq3xE6I5QeqvCZyiw8sn6LBC+QE4hOU0ArYtRWRkZEx4Lw2
08c4y9rCRol4BJb73ogJwxpOCQl73cQSYfskuLrKlIXOrKRrgho7MGOnpD0fPxQLr+9vCJnjzJVr
pNTr1o4nYI9KBOMH6eDntioquJXO0MG/5le/O2vt1fHKWbw0Z7mEJ0WNNTcfuloop7qOohcwrILr
XwB5MFaofTckyxALhETG+xCdpnl0JgEbWDe60AnCBZPWg5j3OUAGr6ao0Vgm+coAd8CVp3LlccBW
oJV2JkQdoIADB2Pbqnoegmj9J9xBeWUABAAtzC81NnzAOYKfyuqo1ESfRNgBQQsCICcirnsC+mi4
FC5wV67BArmmUGkxoWhCwSe9FrbCPXH2l/XbI5uAr0eTDk7fWsrjZhFhaClJ6v//IbvC7FZg4krV
RAUCMRkisS/k1SCYN9HGvDsvcgYIi7SbULV9FCcyuydKMORUQJ/70n0bIcWNBe5lSskb3QmgXF94
txUrDCastP1/+3wNoc+7l3m77oaGgmi30SHXEeycKmbB8gJ1Qlrx4tXtQFmg1Q9RQFKLg1XHRSEJ
Xp4neAT9vQVHDgjAu6MwMIG93R2MqbKd0xSL2n0RBRuiwz9/Rjta5s7yQD9HKfvxU+gEO34f+2bN
0CfB63UWlpLgWvQBSB63iQl/+L+NYAKQX2seI+MrVXpKO5JKUGC3n+jRhrz5DiAXuyxqvbMg68tu
wkXbrmYlrtNfxPgkmkTuZKRh8pZqqz9cw8ZVGdW3529m24kA4FdyvcQPRMvKXGGKn5VoTsDtfCHb
fCeiQQn9MgOMqWQ9KGSFH5WNZYWhr6DCfl5oDBcnw0RYYjlPozJhQ6PunPW4Cf9nJlJaicUaB6I7
SrCcNm4BaO+zC4a12gBmr5d5ULoFVK/9WkqYkbeJdRtENfwWTHbtExBm7dBx13o1q4ar13M9P0Dg
8L+LtAb4WfuWVT+0sxeDuvOUi6gXmOixCNny3nJcmTO0hmomJ2lJ8hRwqTHvotZQG9rGKOUBpQlW
NWrHu9Ylps9Yl2iXQNOv6hEB/zoyCH/+vBTjuennzk6Z9z+FsePKIMxjXAE5FhzW8d7CEi7Z57iV
XBq3IMoqR9ka/vTdaVt47VzZjH1acNUy79+JmaVjyg1dOUw6SlvmxcrYDzTn23AdL+q9zSJGMUFj
DRSYGCrmu407YRQfoxPQf69f1srMAfNo2D3zZMJGEkb3ZxbBGByBiZMPbszLEgnWpa22TurxF7EM
7FhPWuhoEG82AvOqtOrAwacMoncjJQE421iFOAsOSB3lyJvj0uKjexR7q7WDqU4yXaO0Nx8pW0XP
pI6FaHMPe9RmAGP2+jrHCydaysNOdyexp+0OUTTt5ltSttkzCZo3kgaLTW0/jwSem2TjI5XFI3M8
0KOsJ5Z9gn9ch+2rhA2do/3iZACf9XGKZChKjINbg5daveimrTUBCxiMHPguJ+8/K6dcICI+HTE+
XM996k7HhLy6547fLy6oWv3P8uq/y34t9VGe4kIrpGOQZrQHW6338OHnWztW4WKTxZQoldZ8m27D
uODG2sp3PoM8Idv2XI47bStL5Q8lc/tBUNmb/NQc2vC0cH0ZoxSNqsqnE6DNRGm6zm0/KJQZP6qR
Ol2VwbbftMNeXunpXvWZpHej4lHUGuEjypmBehacElTpHrQpHeHxdIHcKnjbvY++v8rDu+t+odTA
tip7IkIYC8eF2F1IW8ziJSiG9k1eHC72lL5uPtUAtDuDJYGBtC1yvOJOLfV+82YShbUmZIo1CGUw
Z8AvuSm0wB01wv0cg0j7cdO4Ey1nJNb9J8Go85aSMFIOGYe+DEPjp6bUeGtNAA5g3pn7qBh03L0V
atkpu+ZRr12ZbtVxXye84Vnq8rprLt5yRYiqITnS0cuHUFNTS/3442Qw0z/tWGhx67O9toaJn1o8
iso2Uple38HVgHVSMZwzg4DuiE9GHcQxOwqZTJwgDYpxPQpegcoDYhZ3O7Y0JZ3+SnY/KKLJdI5x
v+jl2h6mPjsIvusfrY2+nvYd3/wFn02hCUxKqyNZ3fUp+O07ixAeZNAJeLEB7uEs1GcJg7MVztO7
cR8x8M/+f5cEegXTrorYIkzApOhW2HhL8M0A7skn/rUjAP85hC2lAYqXJGyaX1iFGG1rGeD0vipF
0vzQqt8O4wYflb9NLcEsW4hFGolEMIDx1s0lwTjZ4jbysNTo7Mic3W6R95jUVNufpxAhTdAsvoTS
lKnu/q7gJnfgol0h5109eqdT1BuwdgUYd1OakbDpHAT4DiHH4Kk+5spaFJrpiZBHa++nJQWswxb9
+5Sd6YXqPT0nvXXpkMuNwg3mFY3sg50djnOQ6C1zS8eYAIU1g90J+/KfMBDOBiiMC45BSK4euflY
F1pyl1MDvV8tf7w8q5MTJed3FrLLSCpfTos4yBZQDHnIRwoVsHIrktxInaTRFWrDptEkwu2jg3Sh
/btibOGjwb/S8gLSq0Hb+zLj1XuhmoqICqHStZ7jVCTiFXtMcxqqUvgPMcnxaSwnTyOodgxNeR6V
QfYZ51bjzI4ClNGU8WbjHRTv7W/OxV7nGAKg13+kgLliowv1lEHsE2xPm8aZJJ8e1inen+nSXhV6
BXxSuEqlF6MEdCtq9etwTqywNu8c+QQIhy+AQzKBS3PNUTxsaT+8yNcfEgFL+NQJ/zy+wcbCzymf
u4T87fS6Ls8NQ/uIl82dBW/k9cF/Aa+LUqo7OMc9HmWRq1FTFGLP5gbvVzB0RscbVsY43iloh1dm
M8bYydpo7omUy0GBQsI82ib7JJ91fZV/y7G/ativghq2Z0LJGiy3pfHzRcom1ooEJWC86fFUn1eh
PRyeY6GhL50iHRfRA4WYdXQPHgohiDjp02ST/bVuigX7GCcNN9Jn4H2pzvxrByjjFafXPJgXlmhQ
qvv+KjuQTqE2sDkiLKKAUtvSV7BAhPe/VAi80s0h6B7b6Scq8wMSP+B2SgMlVh1RmNd2px4ZS0Jt
V6ROE8hhO0iB/60WiwTNhA8hi5UOq8EX5aBjQb5x9bjyGeECYeqyNejxXsKflz2aFGedZa/g+Ukt
CFGgKfMKjyJpljcA6NuUF3G8gI+Uwp9c0BLK6ipEl1V8tcPaIDEm1sLA9WUxryqPwt9KQmvHDeV+
dx2o9WoiwaOYmIOqFeObq6KK6KM1/rSh+hMNQ7mJ7OFechZdeweApUwNq735+AB3ly8Zo1t4RIOV
prDMNowbMirJ7e9QnzE7ykwFQzxQKW3Ti8HoY8IMfWgRsof1jwfpNJHApY8Q2yF3ay2j7otnE5Zd
Q4neZWC1yuJyOpdusrH6ObefBGm5WFO/3pe6E/VQocRNwMS8Tp5dsUUhc/MJT0XJUd3X6S2m0afO
YRlzqcXvPy6QaMOMtOrLwsUTO5+LVb5JnnDOycnA0AdOkymZ290i28YgRJFRNc2QYNDGgqiBjihY
mC811mb7q+8+MhdejxhipqIiWkXegXy4NDVun9wh6ysnNy3igOrLbBnZqYdVAswmNpWivB1xC1G9
oczo11f2dRV4kUnACXNAbrzR5BxhPx0cAsrkV/bK+mmPZWn9T8kDiXcHuIL4GoDHWfaoeL8E+S9l
rRzr4ZvthPvBuan3q0BQ/kGS0yZAbUPHfep+hNaJ2RHorQazcQqbEtGjX3Km8FWf25P9Ce6ku64t
nGUcaQaOibXvKo9x0qyYtIGg3T9TWoAsHkzBQqkUOHpdCBvxkL4geNFBCKwzRubvF+AUaikFT01R
8ySBjHeiC/qOcsQnn7wGkHXMiXJs0N33rRSnZ72LXM8HQN2+pn5qEIEeikQ4oV/cqtJkuJctG12L
S4pbNQTlLqlrcjp28hgp1hnDGfP5VE0gq0XHrhqHyEJqs0POeWiwbGpWySMLca5fH0WgsCtv4aVn
tMMgQCv6DbET7tuTNjuNOp0B7doFwNFsqN9LjvyLqjBldzq+wJImOF6ZOgk/VOFfsc05msciZ/xy
Fhqjzvw13r/3tA7R0Pzmg5ziFPp7qoaWjBx3DTlwDnjHUssQ0I1FR3t9urvM+GacotG23z/CpHvO
+ObwjTuK+vTKduxjcPUFn6p3IsrgLQL2duyDco4IbhekyaaSyr8r/4TxYxrqpmaZeFURgXfkunO5
w1uYhX+Jnf4dTJlp2neqBr2sNcwGPumbu0f/WwSlEk+U2MACIWtdMRHyAOP+YSEeW3cMpHfypstD
OhFyS6V5kuZ3Pj2e2r9vbEakg7muhccqv4iXaGYPJJ/kbo99bRailD3y03rql6sYkcUCZSFKLGnP
dJG68jWRB83zfNN8RQE+5Shtay2FNvPx3BCeOEhofR1tyQdB/3IrGYYsJ+UadkHapeo5R1JuAYW0
Rr/kHjuHFGqcxl+ySsEBMv4avvE7uvJwEXWDGQ7omKdwNebekTFydBXvtdX4MCFYkUQjd1lzqLDD
fEXNDWMHO9Favl79CdAMzMLRxg4ydewAat6MrUk1/uy3V0XTz6qjvRZK6RP5weYNJDP2wzOjxfxJ
Zbf1pkaEnok4wWtjC1D1AYegOlVS6/p8zbriD6opgRnSsOyv9SA7YZtZ9n+oQe5KK20J2wlsy1NY
Fk5E+hkmB0lR2Dp5EZuFwxaI3WageKn9ERn3F6GeqrG3lAF0e0oTp1eRgJdkVefCI2kV2vCikRwm
lw1JYn37k2OOdYKVWxzi20o9a+lu/kO+5vdkl9utSYRyH5CbhIB5aVejHxgTtNElpOq9am5th1IW
vSGReuYgoGJBku8Wb1tfiEEyQH284bXULHSWXVz6W6ieA5WMBA2OtTav39uJ0ePWevPrVViSMC5k
p97xGUa/SzKIfirlyvaMNCnuzinmXOc/p36kOVNU/lotOKc8VnYKCp+SwYk95y5CR/28VF+zagZF
4TO+tAeKFSxE4sKOvLOqCXsXoRUEkzq29GTEIZ0hBahX+ILmmqtHYWvw2bLqX6KuPodSLUR8pJf7
XS67x7EKj0ORfy6up3x729AUOOFxzo98ThDtOorbIzVCPYyRZe+5HVCAKFyqwA2RJWo7OcVVjqvF
rNp+nWEQuncMapb8+KLG/ZgqmQhzFW0jSgMXlScpbepx5aWtgnoed0WsKphL30lmyKxigSHp7Jg0
SNS+A2PDc+uDKArdL0bhGe8tTN30ZXvAzvni/n324HgOd5GL9pMwYnHi/UW5EVZKFzi9U1WJr/6o
S0jDdiJAIJOLHa2D4b88LENmjO0k3tZ//kVQ+i/V5+EZhpXGI55L4wYXxyn9OeIXhcOzj7xlpEG9
qTM/0kJIUIlWxca0C2xgahDSVgt5gMBxR0MyTNFJ/Hl74LipcmfoM2n8Of8BCCUpMbf6VeQs1VGD
SM8ibRx+8CqZE9j2vTJIsvly6yJCN6r5rKUI3IuCm9eBSwSc/5Y/2zVXN6udFt+nmXa4PP7Q+vSK
IV/dRqWhRySkU2WcPIAcuAiPj0Tfw9xwpCjMbeIBw/qzpHx1ECdo7117SLh0bavEqZWxH4yPIA5L
wTIkBWbAx1iSFQrXOVX4nCAVid4yPj3RCAH21Q69NiZ7jszttlfD/MPoInGB6iWHXa2g4oZZ5bU5
1UWvU7Op2E4ASYZGdBqzg7qCswgkoewRAdNLY/VoRAruOUGnKKZZLPGxb8Vr02aX32hn5IXufkVD
Zd1HbNVvpLOURIUx4U7XJkU2gEysv+8NzXGThuowQchP2/gAw2UGYbMDM2grVsScPdtqs2u30vNw
9IKwq6Md+07JeqVn/fKxgvrfqwdQP5hzfKB5oJCUZ8I8qpOfEFA71pdLdsaCE2eizYGU/vNMjw7y
/qq7DhsdxXSYgU3Lj39RLvZNuWToE5RNwhUmbgJ4A42Ns5xdMvfcoFAfyMVULNbAvPGW4/7laDsS
qnO96sffj25+p0TgzNFts21DL51BzrB/OtTEZZ8igMlIUYIA49caMehVjboVV5coV1FXpqhKA6qt
G4Lo2CunFQDilz6aPI8IrbS6r4Go79PAhqklfgVSIRp67Sea3vVsxwnPbmLBkivLuDuBMQXxFKYG
CKFX8IbmAV0kVan/TZ2nF45d4J/jp8xBDu1VR48e0zvOMy3JVFk5NW7wAqMJ1TXA+jFMHHho2p61
nNhibD6DaVJ9S1h7Lr3+8iQGan6g1Zxzkbi4onZZZvKHxc7fy+5W1Pw1Q3qZ10618AKOx5rmGPbR
pIfh7Rd72eg4EGWW6OY2xflyR0t+n1xtV38lhQqvwCNSo2g0dk+8qeSPZAxTOELPgyDqVYpjEdO5
RFzpmFZYy5lqUI47KNfRZ0+Lp180rE1wsS+kU4EGnKOxWvrZdEq1Q7mmOP2bIAlqivOnTWJg28FN
weqdZANDkYOb4eimK0s+WNnzkh4nLGw/3CtBZdHv/IHAqV/MTH7veCrn2SxZUoosVqToQrkEQqrG
9dE+XeNjCE5g0GIBTHkkG3ZpOuTTSq23ZAqQQpQgG0JC9m19xEicDCln8nwvTFaZvorH7RmEk1JB
Z6K2yYr2TCogH815hvPVPs5LaFQl/I70gVrA9jqW2vul7Pk4a6oW/FVVzazXIj2NqpWqc3luwebW
7QQDSl0mO1kNML/uSLM2Q1Ey0XR0CAmC+EP119zUmjcbC2hOdG8pqevXnWN+FO7/vaGZQ5wnRUcQ
CqnGVV91WB1fwRGcuM+khE43fzje10yUZKvOaABohnndKcQVwEJSAe5eN8uWk09j+9g/W2YVruCo
KOgnTRBxk6lOf5e7uh5RQVZGUxyhXdEMGzdj2rICbvZKI+ZY2V3kC4KeLOpYchEgklHfZ/hfh75E
ECyDcYw9jrE6m5YRpx8uG+TtlzJavDtjtZvlEP7pUQAqAH7MbK20pwQfXtGMhn8iEFkFjQZC8sH5
vq0RYOrrNJi567ynS2Vj7wNpqpWT8I6Ova7NRHkhRGTS0C/mvbAKWzWQ6CNiF2cn70YiWl65Dha0
qphDt0GWz+K/MxWglx0ELLyYGAfWFWOubW96tdtlui5QtyeE5z8jGQviO3nAzlERVQQi9mZdQMhO
nQ83y+OUDt/hYb+zIMsa/3tFAgU8AjDDQFvlIhAhJcEmWOMdx9NrNzE4sPfVslqfKFgxu9jkTWSB
cDfnYkqhNFERtrRvTw50NCe+G3WGywElXFGUXXSRWeivzDcMj9NjPjFW9KjoptDjMpnteYeCHD/X
6Nr6MeiZ7Iy5eWM//Eaj6hRcxigOJSxskxyWedNC5QiG1SrCEuS7RxP/OEDk1D6Z24QPkfzf/HA6
wiif73S1vSQewfqG/ZgZXfbaKqHJlqf/tDkluvjW0CS3UtN/ob19hl89VMrt1ypBzZmnPK6k/Sfn
fYEWU5VzLWxPSRtqrdL8tyQK71w7AztttirnRXxP0tskjdJe/n7dru3wCRPXBpxsJzBsigoPP48B
AtNDoxOmNRxry+YYQzLQHMLUPYQ3W93p/rWHaFxqZudXKDAf2tvEXOjnkQifDXz4zSqR/sgDi8PG
twDC/59RQVikHqSYhn20pmJ2INpQgxDcJ7EwE/VqHEYO2CN+/uWqglJTbSXLogDJ5MZ1ToapoiKu
MwhFtHoTV8tV/vSlaF1zsogGXfHoUMbGhVqZzU6H32rWkOECKYJMqCzWHZQMV0RiieBJYBcE4x1P
kLEgJRYGglhXwx675VqAAm/fcf2uECJj9yIbTRLg+Q2JydBapoIBW9O6HC6jVZWeFmp34oybCFjc
pGE9lg8ye8GKUfIft6AhcjtSa7yqGLuELFLepmiZGl6RK/yQFwt8R7sw3hYD4VKuZeGyZTj1yNhT
TyP47LmoXDnOHHNkkMVPZNYnnB9X4GYsHRc8MXq17LsZ7cNQ502UN2SQ5Qfnj+vYPvypZ+w+WS7c
+EsJCb6mk89HPv15QYlBoZQUQRIB5iFIYIXBoU6buLTCX5Ynghn+s4tXnztljy1qxWt5mSGyvgyh
KC8aF7avjximUBeQi68PfAJ1IvrkYmm5gbv4XQOijgCY2naQ0T54ahdp8OkqZR66WT9Ty9hjZKla
67N71VGgcpC+J1xOHy3utcaoB35/4D8Lv2sTdAMmwuzmVKdN4zSjN0zx67Z6unvGmHrrlOWMZTRY
6CvC05SRckAybNsFpTH7lhN4Iw4UzMtjDyfTkR8tyFBw7/+OQgkpqJX64oVESnJZov1o6vaJAf4A
PApAuelKc2mm7czc2bqHF/Dn2vo8sOiFY0wVzK5IlNDYWxRsoPOOScSRd+y4WQ0lv5bfeMd+1HIx
L8XNcKXX+I2JAIE4UCzpJiDdocciHLtGKOokcujKQ/YNJNRhNfUicIuu3r8xMW+30P2lVQPQrSHZ
GMe0HFJbGbGmJO+DPSbb9FLJauSUNBm8CYWwX7dIsH/ijWPdaBw6IuNVsr+PpdnTlnjCubqXpbjp
hBUb6fjSfuygEnncetlQ8LHKnnU0a8R1NaIS4/OS7WmCbPk80jsNVsqRT+tkm/UcojRu0KIl4UkQ
Z7dORg4y2UD2uzdiQbX9NU/qFkjOxk2C3paTjwhKvca4T2MYNToTQdodSsa5g7jSetD0wSasK2Ho
Ce4940s0ZP7wnE1eydJxA6otjfI1zZaZIJjZpJzNCt5j+8joMhOpvrz1RV4ogVtgoZkay1EbhY4p
4zLA3CL6twzMaxOrPr14sDA9wUNv1GJ+WKw5utwAMpqLek5efpA0zX6EIpxlUWFOtYfVYkuTywvw
iRct0w9hiXWQDtq+HH8cwnf+IDbVjMGbp6QJN1LB/enoaIaDpGrPow8RROSUy+TFkMSc1HZkzidS
03iqaBwXyi2eYx0QLss2SWmJmtZ0Z/Uweg5N9riLQ1qdMqmdPrURBqU39aOEp7QjY4qIh2LMWI/1
nVT7kbaxj53XfCJmI/Bo6sF+KA1FxMyxYWzjrvmS7YohOQaKWdzfI3fRrfW4eGfAtC+RNpdpih2K
HpCAJA/f4z+2ZI6DWYO4JFL65nGrQmlGMtuAzvFHPi7Tsfn0v8ZuAdht2OxGnjiadguULxuLEa+s
MXxW1HV9Lho4tRiMC4cQH/dH2QEVv+pfBqvTjZONGayY1kb54tSU9Z38j5ZzGf+bRBAHOJYgOunh
QYLQ+nGgHRwdgq+VzAy4GZJiJcGd7qgYxEo1cnqKVQiMU9uNIE5rprGm+/6Ucfg4FNH0pyc6eP3E
hH2PoRtqX0nAtchIPnffM43TOZsaLctyFkkEg62CEA0dggelNQ3MDMivcO8JQD/ZcQLLHPPqNU81
pidCxeyCwM9xMYjM5PrWnl3whPcUhrYxPmBmmiUNqgPskakie49EqaLMXYkBgtdPXpIX/imumZW+
odbVZzGp/tlla0ulIpV0h2ptjQZ+jf0T+oFXR9kV7hdAd2lbn7Xp2LT8vIVQf1/ZvuCF/PKx2qYO
TrCavMjpC+t+7oT0vgewd7jlXUht3qnGum6uMWVPcl3k/qeKJzibqPH6uU/03S9AWYaWaw258OI1
pNN+lPCjYR/wTXeUd9rxdJnT8TdVz/fUhZFZaqhnvuBxLQxVgiAz41jj69dBsMcpK4fRXuWJZ+GW
ZvR1I9QNU4fCc1/VDEPZtrry5I8xnSi9FZ0HbgcXXhCJTi0TiLSf/kb5sq0cJ92vi1I/oK7CZU1S
244ZT9lbma8duddBjRu6jBuUbKOquiTPlsLgr5+5kvBduwHJea6vyjFeVlpwW/bK/0sq1uYbnEwZ
U2U8CUgdMccLh2HI5GM5RWCZ1nYdLAVoy46lbW/aKrpfFz7xvKEhvZksempAlHnSx9jrNzuQ3/6H
9XPv+ZuhPsDI+Sb+IxWLKIVgRha9hvd8fPEz/ZuhE91xkmVbedNvecO7coLOI7i+a+OH15H/3u5D
qEZrPMhg8+LwljJhFFD+4kReRgnmwrauIHhA1gTm7SNFLjryHLfxjwS7S6NDY0YlWg8Ky5arzUCl
wtJ3euActcTANLxC8VUTPcRn+VHjhTuxuYnk6mFRZxQKr2cFDlbdL6z93Npwr5ZbXxe4G1bZhGCS
73aeMWOSqSL0dvlocdp2qw/URaksi9K3trPnRj48Z59payq4KcO7uVLjRrG1PH+wfj+4l/rXQZdK
f3m1LlfYf2HXtKMYTxr/+wiRCyJ3XIO0Ap6fpUjiGF0ny0U14Fh/KB7aGm9Q6WOLAYkcgxWD1uF1
9Acid+pYAk1POphz4r67sa2g8L3tQcV9Sb20dXWYC9q6tQ/zle+r92wJMUlX14KuuBEHLdSLS8t3
OUK3nnyv9i3ScXXAIorqlvwrRBEe5ghS1HuX+HJSdDGBfz9zcGavWSehDsZJYosj0stHVsLwLFUr
j02rLt2zwdQnoKpzbTH21fl78y9SZTpmV1X6LwdgvbU+NaMVUemGuiq5VhpqtkmBU0fz5O8wG2E1
rqaVH2Y0RAM/lYF5tQFxkjpPAjiI9Vi0yCd6ItcP8WOSlYk+9cgS0n9sS14prhbicEAlEx7H0isW
VjdqFXb2udrZhcrMwBMs6MjQaVBavMJFkXXIiNJreBQGUMRRtah4W+aoP44IkIudCZJQSsqZ5wPE
uV5ovbrdWN7T9pvC0Bj1GeG2rSzcLNepAbsj7hACCoju8fL5zgoSmQM42NhE8gsIKN/wppNH1uuI
oTKhFlkFuVB0Cw8I21okCz3CwlaHUKSFNL5SwqQEnPzHgn97U5UsbaYjVysiumiLRI4lZXt5HJ54
y4xSBx9Mnto7g84D7p53EDo11HPTgshoh8f4EZJ/ot9ZXHkFQywl4oDe2wpAhZ8cMdQ1H0QVHC6u
wnkU7uPwcR+mH6mjNCO+rQBjaM/lpn68UISlkAECgXU2pEysU32MM83hbq7rjTpeFuWN08C6lRNf
Rc6rJpOBFCudIxn5Y2x07zPog3Q6di/uyMrBFtksZFsNpkquGNhAZ9QH35k3YRRxMfzKRQmW9NP1
/kpseXpzq65zu8uF6vLg6LA2IaRNsWWSOUES/sSttSpA9slPflz+MvPW2X802+ymTAKMWsIj4KRI
iFOnBgEu8HTMy33innRo2peEsbhT/qsqHX7kyTENArPfY5+iGINc4V3hcsOuytHDmurKL3nG85yY
iJB0veaAwfQBetfV6WUJS+ZLH4Aa8ojH9mUi7GRzS5mswSloEK/J6t6Xst0hvq3NvGMRHPyl1rR4
5xBUchQXVfqRTKJqZZOaWRj0AYcif57nmyXIO6Pn+BV+QMLvJR3YGInKroSWelsGhc9EkfR+PDm7
ZVWbwwCFEWdHp4QsibbSE5Vi2ut6nUWd9u/mPLkFQLnO0uLFaZvCmeC6Mvrp2X5RZ/BPbUkYzXLw
TYnQX066cGBaLk2NHAw7WW6R19/CconQRa/EDzL9Vfb7Ps5UoQ3njpGULuY6WAq1vgZ7SDV3nRP7
J5q7BpQLOZ34Iq8Ie/x9IxF/QCg9fzDOwdXjMBtMj45EMY4P+Ht7tTitnhbqOqAtE98x3wX58gR6
vrjPHGnE4xMG/j0unODL0zsSYsRrv76BCxG5nYnIs0IjYVKojFpI2RHFQxTDBXlupiWB3v/UkgAV
mmCkjKUUT/DenHvLTps+SiE/6TVgzaSR87+QNM8DTI+5SfnGkYYpn/+8DQ+3JgRNhTgFbTX7yEm9
Rtr4badRRNIBQGcr1y5AICKBNdpDsTHKM4AlRSBpwHgu1qWIuF82ut19p+d6i31L4uOaFXl8exZx
i8LMI7oUqLrkz9/Xq/e1DYjQNUFO3Jpg3DuxLEmAYAY/pM/I17DBXrpW70hI2p/wKU5GdMvJyDPY
fpwd8dYln3fGxIX29aYKBxRMpRmOc4/SxgSvmYiO6zYl9LMAEKUNEu+unAoe1x6tNIW155OJZiCx
EgOu+k9npCJhQ6CI5/cbm5WksblS+CtCql8DaRFb3TmqL71WlEBReiO4b4/IRC62aIzxOT3mmbAk
jpE6EX0xNQD62A9ZUNTVWbehM6pENn2vacyqlLz+872tzYvyskxCvCWWQ40TcuU2mBA1AH+eP3kB
TW4p7jPRq6kIAVc1XNwumbEkgivzFyUQ0aktUUkcxn5QIsBuoXj2kr7tt+myPpURDVMgYr+q+GXw
x4SYDjtt5/G7GrFxnlvLICpEhwXdxO7o427wblSczZQIraoThR68Kcehi709ou1XK6ba4tpQQLxT
M4Y3NazXG3qmWsL8qKM3LJCNX5o8lSbUC2b+s/t563m1sM+GwKguz3VTbgSwTJuGWW/PwSsef16u
6fYtdZrTppGTvkrgYyeyOjN7wMmmScJRC9mLtV+QfefN57s6f8v6Lnl5u6EnL84OLopFptvurP5o
YPrIEg7hyc1ariAbEzZkJPpF7fk7MOhkBgnOmWaVtC5w8E9kYjdC7LDGC8ntN7ptPArUO8vJ0uJy
chFT61nXL3C341uMcxd0AheIG/pdS0jwHKINAwfznl4wQyGqThAzU1ChVulJifrfeMA+IUd9MybU
BcwODT30ipnjda9hEDOoB2PCk1leZgrOL9GCpMmcUwTjFkHQVaIyfT+HDtXVVvpx5ZILZGybCcxn
/Su1uh/CefbPBl5Qyd1t6LCzYUgv9sOGvzbjUjXfZlBOyA3C8CocLz+Yj+UwlGtRDIteOz/uN4fc
qtY7qCmTCoQgDxRWfLd3EZPibregcM8DK1PGKQ8nAXKlDa/QjS+Or1fTL2uS1w+1SwlHim0Ft44o
gLuGBSFneQRoV0eqizePHjeE4jRi4uRV1c7NHjejICOHBRucrmLbbCrDeA0sKKuQhVK0m9OXDqQJ
XMalIGOkWYQMiXSeCto9ZMI8ktufC/jDo+uqekEw04vnsZfKN++s8fMVo9iPdatqv5OKu2Z3RM7w
m5BfjhEpupVUcrtpliB7BNhSAV9lTKdca2t7gi2tYfSBAcSfX8zU9VBXxZzZ5lU7pBnxrwR/umYY
0oxcV4GPL1NACGlD/JIeIlGcFR20jfI5rogUV0W+Set/Mo1al33hpFkDv5zBpb97eX/GFDde89VE
kEEo6CrBo2VkJJPk6/wySxljS4YOftD+aReinlWUWWcKQRipHrQOqgnAdfwBqY/aVE9doKjevd+p
guNfhX0nIndkSFHbEYns7WNH/IP8YEWsiklnelQohX87qyh3xj+BlYd+FP9x7W1kX6gbRoTzDrvS
96nxvBc6Df8CFCWaeyQhiQ4LgOWP5dt3MaTTlAWQ48uymQ5/IV8U4Q80a08RexEwFaSojfElQoBg
KBA927GkdYx3d8unHsYGwNJDh/pkf+WubqEux5fYfLPapHUQ8lwK7TCj6+fuq+ONnJDxc9FJRn0h
V451Rgpd6dNVSVtOgr3bbpfiozTfnE+YkLR3vV6VwPhrXvMKFF7UuW80YHAZ0JWsPNHBZhQ+Yyfm
s0ShSua5QL+ve6r5iuVg5LbFpgs21ZMpVRa4IkQErOmHUV4hpPhTxjWuURyZqN9HqzKhyGkT8wzN
dgc/vkLd1ZxSfw5cju1IGUM/2up+QgvSP0kXtDzlGt29Zd8K/csBzehc9jRlq8cHFarY0RhyERWJ
NHR4MKuGuBCsm7qbRZikXFRqShYqlp37dyLXAp8uVmpB3zDA3kvNSsv1ttCTbTKP4OU6LtDYUBhN
iKe3ZbIucUU52F7boBvqoWyLDVg66B8TPM4EE6bUgQbjo/bIpM4g0Q/p5zE/JvKZoq8DsvviE6iq
f/d6ukMvlAPrR0PWHwQ8ch85CvsNUJV0I7VOKNfJig7z374b2L9kF3xs91wFl2BK2tGHwr98sEA4
hiSMTDbRmKZ341aEInP8mKEjLwwyJfOPNNr/jAuEvP8wyseSMgHDE71d48jkI3O2njjW77Q4rMD6
CNJfAViorZchOUKnRQ6DMWtAaYzsLYBOURDuixBw/ct/CxP2tiTt5orMlGGr6Ivi+TOP7sI+qH/+
SLrtcInXYTF8VQ8eOXgRLQBWQVSc15YoUo/LVJ5xouqxi/cZWQC7Nvr39wDf5CN3/ydzrR0HdlAG
/RWrnxqMw+dJsFJq22O3iEn58ZMPZ2TumvgaTq1DQvMwKIs2d8TUGyH8o4j/RUgpMM+vRY6bK4xX
Vn6QJeySCnPjwqApr8AWY6H16AM8SaUs/EQIdgJRQ0e6OdjtrHPNKe8AUXYviEZgYMNrQvw0pnGE
lIhRvJDpl7Q3NpW2R04cCRc/lRvEfPYGG3f1tc01XZA4kHtZXX13fs9It6aabtA+a+J2gtxCW4L+
yNk8DiEc9tq7Uz035AOGe6qQb+YNA7vW7Z3FZqhls2uEkW/qwN5TNjnyGPhFcVTibXeEWmAoXSgl
Vjy/4LbV5M/plvOMAdDE0o0uhDf44gsurSLCs7W06IU23uE4xtxxNfRt5dR912J9syNNuElSwf61
MPtWxj13aQioNtet7BYjkLSjKcg/eeWAyO56QOJJ4AQ6R/hQ8ehu9FhdH/11neGGO5AVZKO91PlP
E2ACYTq0zaIto580xaT981Ma6RyD8KbCrgBlB/CDaXGkVajt+KrNerxiKbrrkWzxmt1Af/QsHy2n
M7YXfztnEP96hN294rpOYHzTMVrQIuEmQToyxxLGbI97NAkzqzW0RUQ4XHhcJPaY0M1kbxfoTshp
EJJEV3J4WqEmbwZ11RZ0rymLnCaxA+c8MigJY/KgwwXsXMa3mk8EiD2MTqT2OWvWL2S0RnrjfrYo
fszOO5AdmEfyBnRNpX6fp/v3mVQuYLCuQ9K7vntL4YkwfEiJdqtaoyRLNJPUKnOQvX32e8XmV98k
9rV9zTyn5YKk++h039jyrNx8ToGKEidIOAsqfw82DT1xQeAK9s4fy8Cn7vST3XuCiXT4O7JK0Jkv
4cXyLapUFv8FTNqYKOzlIhFe6VGNPIssWPAlMPshjBIcRWzx84p4OEo0/vpUZKK3j/w6QzcVX9Aw
B23gn7poYWQgKyZWQmnovaBpaISfwB9srgbOu2DF43BRPhV8VnZwG3oE2M+8w/Tww2DX+oPDJHYU
kiLcZF7XoTr6v0pxTSZ1Tpakjq7ONAOneBrf6OwG+SkRoXrwRqmQxc1stLabt6iVqXSNQJrQ7y4Q
VPeLQZ91eiyroSqd8wstY5krNCwF4HlQiFjoUdOMK80f1sm/Iqdik6nM/bmePwg+k4MFasAZVa1W
OtLbK/YqNe2UZe6lwOKLz2D5cPmZ+mKzyt0+GVUIBurthEUsx+64Zd9wtlElc8ZCZzn9WuljIK+e
m9C0qtw9gUwlXoc7F154Vy3qSrVVqUntBE8mtJLOElmKoKzyA67MVw9kygb4mHRLlcLs/lIT8pHx
ATH/R7ttTADMNvV5/I/glq6hhzRgBrgTNT3IlU0XmakyG0TG+GYHQE/U50EJtNUALnS7ZLV6hnt3
eKYICju98cnmaA1Q74Hri0JqQaugWFKy8x4isx9sFNrt+iCgQPBbxVj8qN0cMB3hYksQLj5hHEnc
hCdaBxoq+Djn1yqH5Bt0OgJKI6+qQS/uWNMnmUjrpno//2Hqld38ekNDUDrbDKby3Rdz9FB7La4B
EPhAXrZCetgwxreCWz5cjyHm3v5JAYExWYPzWh/B6d/9hc1NpmmdlgvOyJ74F+XZEVrW7jEHIdZO
ngcJIW5WgsDhKjNnXuGOHDcWvNGAXVuwt5TTadtmfbzm4/tdSbdr/5VRyslYs+vqKk8AYcuKrdZ8
LbxR0rpRsRepcmhaC/jN2KR5oyUUM732hF9l8CdkwakHsvvuSeF7TBxtlGCjIZDzwCy21rjWAzG7
I+o4czmluBmppmNKpsj+HMGmuhKL20YDlnC18cpyrs9tAENY1Q8pCto9ymvTuYwtvGtiiIWKhiVc
WLdvnTihVd+m/KQnNBUXOa0C+zY95La5k+ZlRzptj4gvhs49G4r+uPR9GA0frdgP1VtFj4LAI2cW
hNE+kdo9XL66qpguT6YGHym+SHjS4F8/52xXKt17xJFi5pa6/Af/hq8yXfJP46BgZ3+3g3jFqodo
/Q8cDjJc2Soxn+zUJDgsXUV5HNpHPzKsoKEM1PafrXFkvhnJM66TiR87cqeiBrsr3Ala0IHxbQLv
eQESyeWALklAXPgCOSwI7tF1OOPH5L7soSY9nt/XLsQA7zxk0CQEEw3sO1KrTe8orAFFOK7V8e1J
RGkg6QQkdkxRtZl2x5ww14Q9ksLrNPKq19GqSgoy/eq67iq139rwAFJ6zmGRiGZnvVcIg8WI4EfW
ZjP+thJaata9+SxX/2bhSCzQzcZ+FgpgXSDH+1DHYbCFrD7CEqaKQEs57cMRdfO5w8Bc7U1jM2bD
IUVmCbOM6ueSTEVXA8g+GydEpjz8WD6dChdksdFXi7olXxEFUuu0AUwSnxNSuBslj/18ZxTtmNz9
obg6M5QwsdFnt7Rj78BOu9POBmAlr7px+kLLVa9dnDiuUUD9YPWqqVSJR7wbJivTUg5de6fI/n9s
+avankZDxDDzfxYF0t2V2TwzKMo2Y8U0wJRh2YkVkr7wDgNrE+FHsvgk9cU8ziZhVT+V4zpsIbcV
9HJZ7fGw3XsvMOmHcww/pUSixuYhMSPbXuW8RyRXX1IiSGaGkxN92w0e02N8yEYfyIt/uEq2NmvG
OqoKbjyTBlPQmhdTLhkg0VQ2C0Jccq0TytCjmwWbf6RR5fQfCx4hxb0Sox5Z8Ex6Y1zG3UxV/YTk
yb24g0qsho1/TmOxw4UwXJxo3KbVs6W0mhj8Lms1eaz3gbwR4CcWb5aOz9iU747RGS7E/vMw5fyz
bJS2W++2r7joplUN9PnG20orQCTfnXc0lEjuem9tl+cVqnbkV4tyH8+BLoJtxE3qqN6NmK4F0o57
z2XecWgTvzVBs7D2x9TaDJfkygFhZ2QA1J44QmzeCgI4OSy9JDysSR4U7kllw5H3GvEXUqLO55Ry
h6EnmIpgA0e9PIrQ+q7n0Om0ke6mWG/thwvN+sb7Na8aYi/h1q+1TkqcNZiJAC1mwn3A07dfZ67T
VCZfiuPb8rbKtv4oYaJiJGy+NmUtkPFQ/Ge7Un9BOtxpTHF+d1On5L4+j7TCVAwzRHK+9U7RnbZU
OSasgbA598+6atHDCwzcNxbVnD6vENtBMZuq/t9uVkENMbqdxCp9lmlSF2Cj4NInfu1IO01+Wp+t
839dtQTgdoA2WNC8JfdQvsxAde2XEsT0Pl6rLdca+phOYGMZ4MsdPc+9mn/xVXxoUwpLE0TTb4mC
a65qbTgVxwLgsuUBFlDSxzt3hW4Z+qsBiUdZVqsDaT8MtKYsO9VdcetY5HUDvonYdLaWthGZONdi
8ZsG05MQhub8RQ7ghIvwMu84UamZqTXJCVMdHFsnsrjDkv4LiGGWjtVsHPe9vbA2YrI2acqriwgK
gpVsBv+d47j2u8i70b30yULko4tE32p8AfSCMFlGZNrXa1vEhoIgAa+dWTMyfl+85UiCoxhFQFVH
EVS66Sm2w0e2+063BOU9/G9iXP1wjutSNckfsFZQIP6KReIF3S81XVv/W4Cv5jvciO5hz59ahTX7
eQ0MccK4aMMSbaNQFCmlX1sDidcyh1xoTblqHNX+7HODv9u/h0wL/vJzxSVhLQfX60u30YQRX7qT
fDFiuooYJvsXCx+XFQ0vR7aM1LgS2gwhHuBkbr5wSIsbPSXzLxSHNKKQ8dOI/LnToq3tbLTf8/rG
zkV29SjJC/ZtKaH3dP4maS5j8+roQF3r0M6xw2UrVWMSZddgoOkqODqphBsawPhWSAu+wJltH+fR
KA2MNkMZFehhEyE9Qbh+lgDtWz8Y9z0x7XolsduqbdDDVh4rsYQjHyUg9ctChlEnuz1CRGzsF+GV
WRo1RUJjjv4fP1419ypISw1fQwjt1BGcwNVBot4BvloPlG5RgYvMBj/nqu9h5t2zAfvUo5YjDhJc
qOr7BK4qFkveCCrMUrm2jeAmGi//0pcG3jKtlXzURGTzENVDMLL9TBGJvM15Dr8h/ZpZWfYO4B5s
1HA2gWlnSGDOpH0qGgCsEygZTNAuX4YhxgIpBXlcngDAK9c5kOe87B/vy3sTSWm+IVQhFNKrQ2qk
chx21IL3n1spnmh8bmgI9RBSd0eBZNxNxiF+g0sVPRAjJY9kp/dmV19G4Qp0w9aAqR1QyR52nOor
z03W1iW7Hvyulng6byzIRupUutus8Ax4I5K82nq2Efa7JW5VZJ36W41acnl0qKAJME0oUmF+9Pmp
Nk0La8xdf4m/DNo8StadElqHFOyYKnJwRLXJCaA6NOFL7EySvsGCa9qz/sVoTSX2QQdHa/PFQwfi
sW8DMbxh8vVGfEF69L0NUQYKkBxRISts+Fs5Ygt6UsLQwlo9XzEHQtQAtkKrRAWUnQfbXY0UD2vD
upVOqnCVhg1jmgg+W1MXcmh5Oe35+DdgQUrcmbPPir1E0r8jGovLzQs87gmI2iQwWtf5xgx4q6eW
c6XERy5Qq8qJAjI15iUoK8+xye87BjXXBcr8MDR6W9fFkD4Uq+xC9xUlqH2dNNiWDcUJh6qNuY3r
UIin4D8lq7jpM4a2hvlXfaoXhGaj6AQEMkN2VKeJSWBP8decNI15vcZ9JK8a4aI6CeLOgMnnHw0q
fkXEOgKCEgH+JB3IeVzX1MN6PEam1j9uTeDnbvTiI888056lfJwDSGpK9mwRbEscObdWCMl3sruw
zqLEqYh9qS87b3G6kmJTt9DBXrYJm9L2b8120xjdehqJjCzMKBNXaLyOEM6YlSaXvi7neKGe8pyz
XRW8EyK5dwc5vW0DRl9waL0NynQmwdR5CJcSZAxzy2HIAySh/oZGBjKXRP0oNNkg1yhdFPT/vQFS
vRvAQ76EY5sBEzQnwfEi+D4ha0IAdlDy7Y6SWqOd3LCbHsD42QZHv+zJCWNZoFXkc8LzRCp+UAn8
Hfr8PYAxj8BeGDYk4HQ2v5WAvaDdF/IgsTMU+lX2FpaPJCAshydWK2d0cellopfsJVjbjrGKkcWS
7xJebyHmcMIXxB+t60r24+QpssLvDKXZfqXuuXwNoL4/ozL1kDJOUmQsNDrzqlOjESDNKEOwFuAZ
7BoLCvmxW+BFaeFOPgXZuFxOLzKkEYvDdWG/nk+fJyqPaHSeAkpZU7G5adVadybH6KcCMGTvvnHI
tfn5n0fe5SbWeZrIJ5ueMr+skL9KAZWEdgetuPP6BH3DSUG1gQCN7/mA4MgOlPf4o1Hio+EB51hl
MUvSfTMcMY9iE7kc6spPSlJpREU1FX7KHzUpKwlwIxkCGBl9j7ekGcaO9ccIXtyQOGkuRf8tC9jP
lM3mWCBu7JBchkHlZuosnfN3OSymUa9GEig+XinmEZ/HqYC9lPt/gMM7em+u+q0umaeWSPn4n6xq
ZuS9F4JpzxDImP/c2HHmnyCGwQnjIP4DMVEm7Zbvf+2ZYywVkGBM3qnrjtp60YTRdrxIptkfRpEw
XITmAb4mKqLg8Pe+0IprfBo1a7q1Cpg30K7rMbi54DFJXwfU+BEy/APjXgDBrx22THasc4xeLHFR
WajlUrIJyRKgw1hm6bGdjpeyCRIjVfG5pefgxztauPaukiQF8hnPwvuOn8T+W/SWPW1Jb+mn0FDm
wJn1XcIKHVxhs6MZ5uYWIqPv41uSQOz7liS+9q11DhkOhpdsbFdniwhP/becs98kIUmWyNfV5hgi
FszGu657l6DVQZLJZTUzTs0F3P5jjA37kx9KweAkcuILKBUKxhrxlNV1tkit5DlJGzjX9rezgB7Y
cZp16/K1oiHyxhDsYv1D1j6hfnM/uDkd5wo43urGSH4h+Qrs1EyQEuSDPb1Dd+D0Ub8MEsgeulgD
DJscyiIKaFsQNVnH3kdovAE/WSbN1DA1XZGFfcNPQ3QP8l8s9aIKy7n5Qw1rXoBJZAKQNi+YEilh
if8jpwm/RN0JURsduGILiVHytRJgZ6McclZCkf6G2+Gb3W5+FlEOJwRVUJxL2vhxjW/NjX/Nscna
Yg+ruT3R0p1tFg1dwFylM+ag7cj6PeM6z0AWrUYkH++lDemMJA3+XyscAlK7nWjfjT2tka2VxqqQ
oc2snB0Z1rfDT5Xtxh2Jfqif1iprZzOnCxqjYuYmVHsF589IF4cSMQVWt/ZJDCeJ53eJTk86f7sf
mPjAAUQPPSdNr+/6JKcJUYnALshCBZUKJil/BEQm1Uo1ZfC+GLoz+ISvvec//z/oMa8I9/ldg1r0
SDSgtgWwoRDksSqpSabC5vk0l/0VCuaR2eqeHRYnyMknNnA2Bygoeqe5UhoqqZvXgcl3W9E6Qjxf
TghC2qksH79hlaZqpffKX5DUCc4i8qjlZV1Lo9ThsbBoQAVDvTfjZ/jNHcYvT/Icy0ROB50SHITY
6ZFXJ8E34VGQQyLE2XFTIe9NUdItpD5nop080pDJqEzBeZg3NGTTiKWcatMeX/L4icsntZz0XXJV
HCsZOHcWSXpb2Y1pRoBbkADIwlqT9DBVxXGCXT2iLol8tQuYu13RdInrmKCSiR7j2ln5uLySAPV5
wW762lGsLnbknjJI169m03PtGMbVYJaIfdQx+ug+JDV9vR21j7C0Ceh70oFOL0ErkzcAxaElbtFf
DTwkkvu5C9OM1oEptJ3PfJoLtOqGXRYwa/l+daF/h9fL78kKraJDVbgjpRQxdrh3iM5+0S+bOama
Zk9gBYDjlTcos7oMgTV82OugAxrV5nDR9YzjC4iRl6z7WL+Nlb/uqI3GEUFRPhuCMRN44qEEpCuz
5231cd6OPdop2qFjZFErsF9A5/kOWNELyXFhCawtBMUmPyqsQqQiuDeo9P0YA9u7cQcws8V1pgt0
0v9RX2jFrvY8TscmvYul/ea98BxK2BFRqJszXMHlRale1hDWZtBdMJ8cQA44hMsRiQNo504FhOiD
du64RT2jmaFHtgGIfzewTz16L+zajEKNQjVsXcyM/GTTZZnaIGyy277+jEhFL4lP0nv1PA2bgYgm
y7finnFF6WLxsRKfb7kjf0YP59YbnBQihX96lVXTDAUfDIGv87aif3Kvn5YHRzO/uIrQ2GqFSBAy
tjZch7Q0IIw0eu2MOl18Fn+Yyavxngv3B3ufgItGwcjdPEbT+r988i2RnWapjXFnxMf3TLyTsXI6
dos/U6r5sqK2r+zEfm38tvKXEcab+tdrYtjn52sxT0NM8uYFMNY4Vnh9VNwVsQWz9MJyS52tcX9l
JDkJDZbiSB33q9acC0dUm2HVqCmqfOQ8qA5bVxtl6qqjBRGEsZoeJnNbAXg9GRwumq9YVhpQXy/C
kELVEa73gHcrm7JlaZnszRcWJToTxzgTUwDjiKparxNjE5OkCy4iFlmDhqV/SaNJjxDdFYR0Aht9
gZ8eeLa3S6Efdf032m7zBxIMWIshDTTvWujpCw+eftdRnaVvuUaA7WyWjMtq3RuKqI47MTTR6lXr
tPOaTSxSghZpcrRUTfGYg9Iev4Wa2w1ZHMjXBJJHeF/lOSGg9iFCzbq6KyPsSKOTXSgrevIoDpLE
Pf3VibNdQckymLuPNDEExXWm5fFito2RaW9Sd5P54vGXyOPxRxVI6UHTYf3SpvhW4B3h8SRfj8At
1ZpzAt+8/X31y/DH5kRU6VtQ0hMK8VKnhPABY9aFdGjxMiVv5tgx+3c4BUvdXYYdawiLmfY3d1Cm
ArFwP/FCDIXSLd4+UFdZxbV9fcahonNbEOr6DyfEHBA03FgksfWpTw++0/8jLE877p1QgYnF18bF
VnYtjVShuaymQWGY4blA8+3KnuNAVV/94PB6dsBX95a2PJQ+sUc78P5NJCD/M+/lEyjhaVztmJr8
8yh4ph0qtpFLm1+V/Oa8hHd1jUCAhsi7jUedAIhLKGk9J7qfA8rc5LInbHKiLVWVsS9ywRJ6SWZI
QXTbl215R3gX8+/uf+txB+5peI5gamBRC1rulBcbKL+w4cZxBjrwQMfSFXgrtzzkR0HIkxCf0NrU
HJMbARyUWSS0N+wZlT7yh+ii+ks/fH4qJCpzVmkP7cfOtbnnq3rTxVbbgn32EaIjYJKz9jTvcnHC
q6SRuW5lKv06kpI1LegItsAieaKMEV0He3AwTa1HV0hsV/hcRHOcLTIGsRWacXEB5AyXo/P4vgfN
hcjXlVL7kcKNfNrgSQUzWCNo2AVjrHU/FGd+KmAmeo/+XAuKJj2VQ7LcK5HGjMIoiflho45ZezvR
2Nr79h7ZWsZTA+XHwM2nwW4mYzVxEPArcVhM/S2teiN3LHe0nnPqRq1oLvg968F2H7VJM7bRj4zP
A1eG4zyIOM7gFO0dUjXJ3Yz1PAuJMPsdsnLWSJuFKNaO1n3o7LRiSo3lltv7bCaJV0s1jfgxb9Qw
c/AkXURjlZUu1SjXIj9msIxwnfICnhMPw8QRFh+EaGQej592qS2cwodYEFXHLqtsKRuVKmazVt3y
G241Mp10q+/e3r0zbbFTYeHSZ7ymyaOZGa1/2hK4TWnXz5I9aOscfJi4f9mW8ZYsdLXvZ+Nb1Whz
BN2XIFRiWSiNAssD+TlAw5VsiUv0t/m5kPZQk0KRde9cvYP9eNyTov3fC4jQgiZgCCn3LW2Z5/1g
pdQpRGBYSLmGXjHApna15oz5o+NMmW5PaBLyd5naIdtTDRRda7Z5LP/w212jUYYrJZTzjJnDkMLU
bjppIOFR3OX7+wP8Ge/uNc41XuTt3SPJ7qrUST1cHHMqVoau8BvctngZ77OoNpFwCVmByIvzhBQE
5qbfJGGquVvPUrijOmSD3ecG4VYVbcGxVozyWNEJetl9NY7Oh+pHyXlBoubo1Yc6ooiJYcr96AZD
MtjIbXUXaVLhFnxXBMD1E9HxwnpycKn+A+bnM3E+iQWZam1fOrpm9YaIh7UMnU54xW/f+qiCM0Pw
aDHxP3Tm22UVQyJ8J2+F8Y4rLp48HL/jrsu0oVWOeLfS55CKlK41LucYYUBOAYvFmcvP1dXjAk87
u780HI/uPSk/h2ozRrC4AdHhX0fcMxUdwsdCX2zfaR6kBLVoD8rbq6qtMUYcCA15zN7aBsBnGpWy
ndX5nTqAz7u65E8+FY81xSbWsU+RITCowFvFgtTufrIaxHJTTbmrfbNNG+LVGid3Ia4pEd/KXZr7
EzgALTowyn/wGJr5oyFKgzUSqItInlU3pL2kZbzVDqPolmkgiPYmolj67KEXP0W56JeGxMoNj4lq
bOr5m96p2lEkAidvkakwDSeu9NOWKDVqUu51MhJBt6H9nIGUFo2S//T7K6AbQi/ojPzETrI5clsr
bpkL72AmZZ3dkX5PW8xywd9mZiYlUZvIpglseFv3jFkiIykm59upqGr3HD8i+zBqKiVv3tEn6Z4N
wGj54ZQg4RV887DpRdPALshMpcOXV8NCCeSPh9j4Dlek2wKPg55tY9Ym9fOttrDXVCZCWzKSPH9v
Z0UdsfNfhSYqJkW8IBn+cGjEt2sXvz94ZxszDHM3B1Y6+vSGPesr7WUUb2BDdR2Y6kU9t8dMqMYN
VRwVKQBQFWDz3vEUuls1UDEKZPi4pUjEhET3lwCYgAkGae+6tn8Q/wYe3EAuZJvO5oYOFyRPOFV9
K1Coc6pzzJE5HsPu8H8jdXrm7C1a2VzEdIrEzT4l4pYzv3JDsUDU0nvLlGVm2oEjsPptLd5roS71
/P9K6nvkRg0Wr/yXgYku1WW+N3rDCfFeJciwmPygPCKSkJusoczhFfaq+AZjcjqRh3PgRcUwi2ip
qePFOIE5aY9+gD4eqFs8f3PIQOB8ij+5aKi7UkVblbHmry670mtf7mlNrO1JNSF0LAbEtcmItDav
5EMZYKTi1qokyULZbopwPC/uPL+WJAQRJBP8D38yE9get3hIcdBG1QhPbZCmnvA0DWC8HG2IifmO
tPhcSs1umUpyKRcBj9IGuQUVUcxCYUJzulPoJp7LBy/4i+QCRzJkiYxVRe/UipIbBqTxen3Z8L5T
w0J1Ij2E3KYsRd+PqY3kYSM7cPb9OVpc5IcPp0zU/Pun6kinGESZfMoqWdOBYHhtsJV9FHlKLcVR
74Tiqr0B3bvFlxklkEdncJebQGsAeO1A9HuDqIRPjoalwE2dfphashdKLP+2NNA0Tva736aQ6RIN
wFBznLU5Is/z6ESlSZgnBH+E0zgr71RnJvPSJGOsa+6+XLZpOsXQh00nzyfqD9qG7IVhYVzDKl0E
yNTbXBeWWr+5Dyu2RJhqxtNgqnP6JNcaot75jB8qecP5fok1mOKCckzb9Mf8xW7n4lEzWDF9/d4m
acMD/Ty7/dCJYrHcvOsTjlTo9Zu8IDMUJJUWECfK5JEt3qY34BFLfnHZMtZmJ0ZTK/Gh8KEfbUv7
i9DjDqBsipzlWqzB/lPdRbal2jokQbhoab2aeKdFCCMWXkBsW5MT8/F6E+RiSaPEPKoJ5T6Mgoh2
pR4B5cBcg+0hICz8q9dzRdOVXXYMCp/wLGSzj7pyXFtE9aKC/VqZXRhGgicRBwGMGn/7P9qKR24H
z31oFr3zajsdcqMMLEu/p5ADHIuyb0o6ON2NqrxU204PlA3JcHN63cBgA/5ae6TV4kpB4WYRIYph
DL70eiw0Jx0V3pVmz4MIzg8v21jOB5f11DdXJd3XUbwOPEkKStckQ3hbOR5PNwwzM7OYg4LleMcQ
3NU3JC9Pkd4f9oXXH2yLb0mCxNbvHzDXEU+a0CqnoIBfYE70ydQzLTkz8JagZaArWQrxGmqaasuO
c04ZnLeNPBX2BjB2dUWcjrF1C6JMasUhG45/q778WAwl/SppWWNOQwWN5wWvREcd21HMEOwedCFJ
3B9IFaeQ0xFs/ZpFJcMZI4rSsvxB4BJk4ejG1S6WpPEllOM1TUcY03vyTOlqPBqnHNdx9jbs7cXS
8447pge4kvQDldnRObaEHD5/TefbgvRcKJWs4BHTHJLgF0DIeCMIyDg2CB9rlgacl9YZQ0BVS9oG
LjcbkK5aLZfEC+825kxtAmf6MxVBVDVxugxcNbz93XCfcKX1CGUmQ73Nw9kX3/FT/5B+EYXrB3BU
rGdP3kbsh//pgZgxuIoANL4Lbw40Owhdy7ei/lY1Z+EDzo2w4trT/ypouiSBMPWqXqYS37TE4qKE
3fzbMW6H0PuMjLob4B1oVZDiQdi81rIcHtWLUNu/JZnwWVU3zmN38+NgLu6yI84fMOwa205zPIsw
o6wJ9+LfSIRrKUxsts5Dsz0ZhMWwRim3s4k91Gd02c07RkojrbtCTcz7cYaun7QlIEutccTtfneW
0+5m06D0PVOMVLAdKZxNYRgvaEpS7BwwkAD7y00ITocn3SPs1G0ud6ZImcG+mpZmczE1lPJgjUMD
YwG9SIjlzewFYsft184lLg2mg3Pu/RCDeLwyfc2V3goC0hz2TzYilRv05SI/CgP4/iyUgd3fkJed
EDL8Zqq3Fx8rPqZR6u6m+CQnQjk9XmvdEoYB0Px7OpJN5X5KJaJyBqWNAM11uja6rH2W0QKOJJ5k
D/8SdIW/4yzP4hXUDnljodGUqTb3SLl9IXVkbUFmVGO8kS5SQ03EeS3EGnEwZ9vnMxdup0vCrVIf
u1nKpf2sohj7vXH5sLLU1G/UnZWy2jELnST1cu48dRpzwrpT61hJUyNOpECpK3nkfaTKtI7NCdpl
Z9jUyWaLv9cXYoFwuY/3Z3Hl0Pzyw2v4GixZlFNUSqBgzJOsWV5/L7ySWNsJVM2GcDTKfOL/eV1G
FiaBNdXwodBxzxt+feuQsJMGvUdbW1fU651C63ToLLe9x7LDzJf/YTwKLLFJwTrMOYXLpdAC1r4g
ztPODFMa2AWRfHf9T+n0NU23E41fmE2xLmPY9uiOH2jBtauftv9HxLpDWbSt9t+vr50uoXwVg5N/
vxMp79reBK1ik3F5mSy4Vk+ZTieNRcjwY3iiuUPMejymzQY4a1rNNgpFv9cJs7yoc3gd5KQgfmH4
kMaPgKAebg7zJmSscwjhlpfptgs36Gpge0JyNgnT8dvQmxXXwZmWe/bLauz6HpM1fXjif7v+BWSV
H6hKzffOsLXXbvRePGuSyEeY2B2S7xHR5KMFRHSfy6nFcdXpk7BYXqNMdlyKuJGutMjsjRPlIOHw
AEi5bt1BlSuHUz8Nywm7oAyFpLzWTuLtray0Vv75LVz+rek54PSKtgLOlknBwc/zEO2qTlT/0yhh
SxKwRM6OrDcH0HNLEou19aMzRSQN8GV9OfRvgX8GefDXZZLBMdG5U8SRh3ji1a6YyUZDKkQ3MJT4
mchw3u1Ir9oyylTiH0jShAAeXdG2nb5V/FHzhyX7F44DX3Jqqqe03yjiavAS1dW1AmsCaqg/sFKK
Im/O3cCtv0Bf9H9diDWZqHt3mdb2P/B72aLD85mmZ5KqvrZrKGLN5ts3YgEKIYZpMK4eYpRfl+nT
sJ93r5uAOptdmfaHKfI49wa0Yv0pnzGSlrStS553TCbY+D/CKOlqhqfgQwxlhezxaZQ097pLaInx
UdIWa3Xf8uoW2vAQIrqu9Oo4Imupg5Z5s6E3wYxagreQSLekuSJrxfWSn5I+Jd15n9WY19ZK6Pmn
JqHDiZoZ3RsxAb7VHGa7w2JwpGh7kmDLhnmXvjg+d461sewvVIQ+kmyPQA5SdeNy2dFg0ztcdrVB
zNF6c8rhjQjtoZvoBbs3UeFG4eCS1sfnjz2bRhvPpwmC7iXzgDRT+1egPeULquZyho/JGby6G8Ca
730jzRq7u8LqA1cCxajUTRyk4SJkJymmAW6dIUj8zY9xgGaIHktSrelcfK+ew51KeSi+WMkUceC4
b9JylIdHs3dBjNK9i2Bp/apxTfcEmCEjUYMWTLlvSMcKRTERyqHSij6/Yr/Lk5YisLb7QzMKy1bG
iPBD0l04xRjGG1QhmJPErITxNkmf3j5BxWl4s+zjFvh1Z04rgTWYtL5U3BYnh2Je5kd9k3ssQKjV
RMtOMA3oA7lv0Y/Mqxj6JoggDR4zqD8gO/Rh08EBmQ9vboJwLlVQo8VtP4gEWnU7YO5FHYiz4b4/
4JH1BGDfh4Fww1cPDh3Ue5UzAUX41FftzpdEsDbVGEUUcL+70/L5GXa3HKbkdeEYfwduIdsNxjQ4
pISUCSvxGeaflEpM/DPSRPMtfxomVFV0TPABqWrqpsfTSLAggKqNWThK+9LYccCNyorL7YnGwD4M
6j3wbgWNy2HoTd0qDrUgFqkUkRYWzJllTFf0pTBl6IV5SjlBRuLb7KDmQpITGbDkcvnvC4HIh5pO
eAT5olhzbfysLC1v8oAYza9j01smxI4ZU8YyHd3Tjxcw6k6bFC4XvvQsYrrrKAypC41XEB7utRYb
Uj8pWHT3ydZSXkA1VmULIIt3IqEglzA3ZeGqC18cb/V2FNJFN9WB6orNKlbCq8cKvkJFsQ9Y+BJ1
lXitox6uZJVA6Wb3Zx/A49ThPQDcw1UE3Yu1JmKLxr+gszX94XaRliZzLQ5qBX2Wkn0Lq4Hq5tRd
YwiXVu0Kjqugvq3BoUypCZMhIOVyKozm67qHCNXAsu4iu3jatMgPW/Lcyj5m+/b+u7AMS9VjTpW5
UKamTXdYLA6BU8Tci7MHYi/0fw/scygWuFk/FFHvjA45kZy1UVKtEzXH6SnSZsQSNYlmS6SOgwB7
Y+3e78erDOLOWK7Z9EEE3bzWJFBG9uw9+4uY0kkAE2hY6gXilkvRASIP33ebDkNoWKGY2utwXudG
71QKNitJ3F36++dh2h7f/ZPZbJQaN46VnoNlofgcBZOaKwAy/BQhHY4v0wJcbMT8XD5XQBKrCZw3
osRd05O2MC1slneoqabMhkc4XJCxLMSxkecCrIbX1Dr2OXDj6UHHS8ePNNwiEk5T5sU7In/26dK5
mK4PTaV9rPiqq/1kDsNeKWsC2lQBKCCYGkWfiSLz9K7WLz0aczU1vGeUL4tPFgPKOxu+/b4P+qkj
UzmYj3CU9q8sKkwfyNvsX5ZxJxRgYJ6K2gKa4GAlMQetZMu6+gf+gL+brKFDQw9ulhnaFKLffWvc
t9RRnr3/XWDWoHEwcQn8gCf96RvoMWCvphAijqoptGJu2HHeKCD5uP6Sg2h4DtZUHY7xtqO8hNTk
/W6t0cnOp7Lv59v/Ht3ZFTUawkjx8egUyuu9GJO7necVhZAkWyt6x5kGUsphb95+Zv6u6c7AcwXi
JABCBz2IRZFXkhItVNF8Gn+CNZiKmat63nbbkXq8QRuuCsRAavXUMj5QrWeqPNmMRu4uBe30v/DA
mC84N+7RuJ701yCAi4ZuqVd0Wa1Ft5Usf9vUXLiA7nlmUpRJrbRfJcK5oxS9tDbWfvkpCAS0n987
BWcO+94bM830leRPK9SDOkxHvgbhZ3YuNTKwrm3OIZEJvQGMO961OOQo8MJMTZ31S37QfviYsFMF
bqSF31k3gBSr2KajPvbdhsVzwrF7sZMwGvzYQmolHntDCpifqSHGy5Rprjukn34iRxPMMqgAumTo
ertaxT3qVZ9cN51hLqgXcymxs+RfoMt5rxk3J0ILC6BuD4es2C0UhqOSzK/dpfF73rOgNK0Gc7Es
AKBcTCAvLJyKQwMtVY+GsPHbdzPyQ3JdLaAM0yEGcByp1ERejHgtWb64UCPkGRf+tndvztbrTdKI
5p/VWPjnaNbqvB+30C+XqzrR+xs6GtKbsNdnKSaRm4mhHcwxS8zEsfc7ixOvcOjhdoyPjte07yAE
15gcejhu+ZD4mdXpj+hMyWq/LGQtqU8WsmNgzflhx9xNovP9dj1J3m2cN7IQnv5IWxZYW+ibMU9f
CPNT9ziOcfh/lLdShuzPSRG6+fUYCf8CD8z72tlmfsdjney3AeLGHfunRzwbPousS757FzQZWOdz
rpwdjVBC1odVUBI7cvwzNRk6C9+PMWcNG0yNK5k4GQaFrfWkZOVmzUlLIZJ7S3OxrFp0JUvzq8fN
xgSrC60reUWOc85WaXCHfFFfjTz1GkPhdzwSUKekox2qwxyprYrws+1nYesB/UaElefTiMFipqNL
AnCX2beXeMC8WFMwGnrD6pqS9uN3YeMQLhSx/8pIUfkY+3gZIpg8GNI8sV9Wa+4mzQ0CV3nFv3O5
O0wTWTJeueoEU6tOVeR0mobmiGT6zUHsaozTStSVR3FEMNy2ojVdXBugnTMvu9U6+8/2Qn7Df3np
NxQBV0LarJ4GsPSwHR9+LZvYMrN6gptUIgfFz0gRd0utKAnaDEaYerhYQMHj2TKRjvyCq0RoyQi0
y2hio61P5WYqBhPhaaJKY033ejwTEXOF9OWieFVFlO9K1vTZVw09RYaJIgaYk1wfdREsvuBqhl8U
nXE8+Mgi+ja5hRYnKlWRO/l8rSvdD6v1ltxH/kYor79MxJUSQOw8XefV7UEW8QgE5c0nfQv5MGd8
8U2nSxBpEXHhPPQdQmbtBMUYmrxyDXz6V2V20L5uqEfYuCA1c+cHPb/Kdf3Dip4SoRu4HZl5o6oG
11gLrIknCzCzWeJ5jmLgkZmS95kyyU23PGprOPaQehT/taEBemY5SEHNUSLQT2VepyNjJKa5mMGB
9RutxtJSn9iCzbcZOXilhfsP5DOxHLxJi22jgbBM1KsD5C/eT9Or+EUxfvo9FCr2sE/JXml2Uumk
caA1IwHlq8qwmP35fXHAIx5jRnnbUWMvT/vA9K1IsCHOvScTL9Luc1DhAQUjeJtRdpdGfJFqNC9K
ujqlgN4sYyZIvGEAxpmS/6l1JPucgc9Ongm9SoEbWxq/cmAzsQEMhlauxZ0DHqPoaq2wee/XpE6q
MTdkL23quXDjaXvbxWcRl/oGF2aB9YrYOZA+bZSLDJf/29468FXfWaIVu5NG7vTuhcntv/X+GcCQ
zrzZ+quu/oIY8J/kPbg7DhXAVeu/JCnmvGGSVqjgtqrTxbuoaBPmn7pu547XzgI1f2Zedr1wN1Ma
idIvspK+GM4arLAX4xZxLGAzZVwU5fEGmxKHET6cMG1rnGy3MXJ3aCETiiQPTz0lzaMegzveakvu
xcoUuju/qW4jgw8jF9ki4e60IqxFEI1/FXyaTiEX3G1KodT+cdO9iCC0K6C88NfVagPvnWeejrxc
aAqSX2NOhLD29qPTbZGiqlpw6Cv6JTA9+/eC0TABmEDDwFJh0eFIOOdjyPZfYUzj1Sfh+F3RyeQs
NitStBaMfL9vyB4aSjBHqfEflaaUKGMzdIwX8gzwbeDjw+Vs16iAfMqbL7IxHrC0l53gHkYGxn5/
GeLa9FgASy+26Jh5xZ4Z510077qR7/mFWXp1ce3+GT8h7UfuJYtSzoW8qm/qpld9BmpBCdESqYHc
Fft1UmQV2EuzmPVBiw6g9k4XqGgJ/it0ufgxDwv+fSh7oKaX+HBhKo/bYRailFDKPc0cWb9Pza0m
viu4qTtMthLDFwGlWazk9NdN/LLbMZo7ux+oIBYU19EYMS+hVIAaLXIvnUAp2RcfRtrvcahjbuvG
yFsQhZFDo81Wrd2tgJeapaEGB8KxpgVEwApPZMoEnrjQ8lXsLgkOzkDo1sKj3ReW4JEMnbm8UjQV
D3AEEaGr/h8gaPWJGAl8dVzce6x8SuUFGg12R3ZZNCFMu0eVSPQPngHBR9ZteMsaFAI9//4DfBAi
3ARsUdiLBOVg/OyZyxn/KZuJEYzCc2pc4UoLTcIcJrnA1pxbI8YjSy17+yiwpZU4G9+oGJQvc/d0
e0OzgpHApBQNafikq071f1TGGDtA2th6xgX/SiASiWqHmGIKSZIteOHs0hnIF04UctTyyztLUDR9
8SxXjEdrdszFVTuyqhbkSgNHYJHwY99vK6Ry7vVx5KHpQE2Vbqk1c6zjDmRd2qj16KQ//lHvzrus
J1+lyEeOcbaKDg1fg1IycQMVhVuA4n0TtMtWJf11lld9CkqyBBwF+kZ5KHXl0qGVrd0CuznX9k6R
HI961fk5GLa90Hu3xRdgN3Sf2LUMgo5ykCRLzhiR0iWX8bWIDHTJ050bIFA0XQM/Ws9T5+tR+mAf
UtAJqI7of6d6g9oGjsU0SUcoITDjuEieTA0K8Z5D/BZoB/q4AO6ExKB9FiJgOICa2s31QMtVAill
tYXDOR7N8wAS/MAu2InnktmmAguByx6gB48oHAbECU2iIzcJRBKL+6NlorecnKv25Bklpkjy930M
G8Jh9QiQDfl3Ju6b/zM3Ymvo+/WD/LXT1uKgw0ZB/qpl6U+s1xFg2MQjZiDFx7s3/nAtnZfzEitx
1a1rBWyOrSd85MY4SpZwCtbozO9o7+QpaIduH2vY4/tjiHbn0/1JmEfo1y2hcq1r32ISdCb/eIJW
q+WX+4t/dfFelU7i3X9AEomKhyS/usNL9DsbStWO0LIdlbG718WnQWKuXEKG0qssw5pUtdq1G4Dj
ZzpdjXKcMZKVpxx9jdpiSRsbqP40FP67+hxdwu67s6vw66lQMn/pncLPC6XLjqCtxkkus1xmtdy4
NllhPvKeBIzbDUCb9/+3G8fJSIaJkXoTZo+Rq7X2OP2tU9ZiGkI5R+VxoUvQ1dsbdNoIqKyG7+wZ
jFMj3kKM+MD4krXrsPgzOqQalPJeOObuxQYWWtD0aEL2jvHRs1aH9vv9wQ2L7462ayzESSKlbskv
8hVCW38uCW/0kI1fJi5B2WotBKh/IjTQlOWCZ8b8X2vYhFBghbFGI6a8G33ij+lURRQdUcgLeaZl
jgy7EiBdinIHpZOugzCtClOulGn6cjiTC1uAzErIckBorGm0Id03eXdMYTP1WC90Nt+GZBA+62te
ozA1wHu+L6KQXAv3bj5hm4zDucG6rdfCYcLitkZ8YFPwDO+/ig8jJUwua+Eyv2v8GuXRUU9Y/MrT
fHPa0LdN3Yo3BVhN5HKwFdgI2iC5i/SE4Jp5ykIYgtsrvM4W8BDY9ibE4iN3aU29cW0OqIb+qwDo
OhNBJ/nO7+8N69B4ATC+TcUPZwVnLRXnNRkGjQPjNxW2PBJqnZWeOXvM3ZoZVBCsiljhkjmWLN3m
bSZbrQfIdwqPtdidxGKWL5z8zTNxcKF/s1Iq7wSJpiJt/uKyODgPMMFjQsUVrDgis6baivXPw+dc
Y2+STk8bGDBw3J7xdUXjQbMLOutS5ztRfi2lO6kMPeHtlnNR/P0tOvWCn5fi3kzqiJXqtAt+9ds1
B4h1XdHWknbm0MgoTUCh1uknGUn3vmG5g0nrkl2rn2HivzpPwDDCF99lhyV4E7eXPXPCR5XKhggQ
Y52G0zVa05LuXSRMD5yht8Mw3LrqkCTpc2hey8TuRLEPGvTZn51v0gmdJVu8fneRhbYWejFJa1tp
WGDQYXuhTQ0iwMuQcKJLwxhm1RdMc5HyOenuDTS5Zlmm5yfXwHGPOG8KOlVpUawI8tHVpMfSZAiU
Bk8jly3Fy+cyngM0dDLeDX8HzRfP709N8e+L6WSYSBFEeyX2fruJ6Px8r2I4fqJzqsg4SAOi5+gE
DOsVWToMOA4/S/vxUL6FktRyfcWNRo48QxSwPr0y+vDXSGkfap/ILcKONMM9++AchJfvKAHbtcyO
MPk6/OKf2nzL5AwvH4EWEw9lwr3XysoDEKTtXEHTVFl1YpHkVFH/x4XUqhJ453p1JuCc13F16t9R
O+OjdpYA7PYYfE2SiD0LxoncdoSDLgLikRcg0ARTVFHRz0fBK6DwqW9ozJB4SOg54zA/Ck08V0oF
jaYmtNY/VVfOn/AXgdkmn0lNJa7VVtMNQMCYJl039JQvg3HrDqqD7lGFnKou1mCbyQv2i4qsUMaa
NAGkMW7lIg/RP4tJmg1O3pMwzqD80k4zCJTrKeN+NeRGPzhBG1o/Js7z74NjsS9dEmV+ejlz1xbw
82FRjqHHdXPSotYcpGgXEbtACH971IrK2jxkO5XKP/TO7pN+7fPxhPiXZE8wynN/J9EyXmVtPAMt
mPWpjqU8e/qGFLJJXNRRP6gxRqiMnCjMlCE0PZcx9oRfLVzK8Za9DQrQ61TMLWfN17GO1juSGMJh
Zt8pENvMw5vYNAOu67RMBkc7QOEYZJ9b39F2XLMR0/auddvsGWpFL19LAjQhKNx4ztFnCgqstfCO
xB6OMrxuahwoNr/mZanvQMBu69HKcWJ+yB/AAvgtWe0WX0eqgoxnMIieGWtMofshC+5KXs1BJ1vk
5nNa3eZTMcGjxjGQllIXhw+GA74UKxGWxY1AHx8UefTgS6ulk5EbglVBKLV/kWj2btbASXniWMQi
4PsYhKsIVNOXYdxInU0pH9vuKWYwZHuqHKm+40mBmBtq9n33oUknSdH8IvPrV/lSNZfsDN9fQRyS
2a49l7SDhQEyjX1KhiRLtzKhhA1Q7w3+XwourcAJnVtNJ3svWqTqTKCXJFx4XCsT+p8zIhPgqXbZ
QJCVoWTvgiXlMnG7qAN+Cexv6Z0qJmlp5z1mu/VLFDe+WdoB4hoeZU75szrHXx15h20/qt2HH9ZX
jxLYrl0bxlxDThRxp8xxgvPdtrgNqXSKKmYj9uSGgvJkpcl3CFFXlxuYNVaF3QvOJdijYONCiugr
t8es4ekBStNXE3tq1If7Tx8Wx9HyKumx5i9W7bqolOr3QBS8lIBaFb3TiF2bfhvCcv4hvfC19ELF
5ddVdn6EE91rWIeSgEE2xhnM/vNHQikx7nr8kfM1Ejs+rCBi8r2gI6uWeglI5fh7RCEvsd5LdwjK
QpappS0l9k4lSOdWEP4sQpqBPQkxcJtXbsU5TxxJjfuPrsDGpThf0CGj0p5xNpJ6AGjDtRdfHzte
YnFrqqX4epep3LwYHdjhwavjetZvJvi1LChgI3h5HSFV+5LDz3hLzAi2dh5d+6juI7v56N2YPRPY
s6CsaZIaAxNKdEhateuxm7AVh/hN6TlmSQqaCoJSyxibhHIVEcQoygZGo+zD6Mnqxz+KAxc09GEG
2l+Y1+rMOpnNvHZVT7KJsQk/gGgQs1k3aKKaX5gtrb7PVAKBGkV2ecX6+/1PiEtdAd1vXkYDgoUL
yqlZjQ0Gdrw75V5a1P0pIuLa6gDQ2dgPQZakzkIu0eEEyG2A1TUYXCMROAzRBQfJMdI2apicgt71
XYZJmIOIYe+h+i6Zr9iSHWb+pj6I9LB3CnmqHoRTV2gS1c1G++AC5vfRkTNhhpDGmypVnX2iN2cE
mn0bTRtphb3AYoBpleBscGDvMZb1aeIccPXd/H0fNXTY9THa6728EIztzpr/rhCe3W5v3I/w6rNw
/DIXGABG2ql3a3VxJl19RzeDqr9HlirLVPfxzO2fgqV+8+RFsnpujppR/5eVxfDRQbm90a9G5NmU
eVodKyKj3jKHdRxSJx5pUyyoLbUnu+VAAowME4EOB3YOSwSt7OGe4M0YLRCnuo88qp0WR0HKz7aQ
fKy/JrtK5YXgt98wuUdHDibLLf3ynvFeMDIthyknbL4UexJqytLc26lVLzElrohfmcCXZiAjSpbY
flMgSTWhp1WLtcBUtAh99fkMaoKEOfX8cM/3DMDJv2YTgGukCsLMkn3KM3aIQ0CD9nH2PxK2kV9Q
9nv6TnxTypIrm5keucNOWAKKtYgHd1jiB2eSoE1jqeFpjp9PfUvrstFrkBhITOz+GUMY/hEw1zCb
TqPktPXq0FO6W6XC9as9Ddej1ASpC0j2BMtve5e1fc/U0fuzvRsFgOdLiIH7+5z5wuu5vpKGXy5K
6XF8voxTZYrz1qgggof3w/AeKwPb6+WSM9Ra9o7IYaaNoQ/dTyQTphPuH0eBYiC45wCK59nw7s58
PCn3wi6c2dwex1+Z7u2RImJ48pd7H2mDou0sdigLOP38UjannF649mmAMjxKNh+a6/eoxp+BV0fs
9fRQVN89EU4Q+2UpTfgtwX5VehzrBtozYZeH20eYGG62OZPhiG62Z4xOIfkJ51FeJ5wNwp3UKQmp
8PF4Rp1jTJa/IEFc8mNIhuyAxWfSOthlgvnYUbsexpFQzayYVUD/TpDjucsLu4BTtZoDYCoFRmWE
7C8luYbBk/QlXPvD26DdBHtPrIc5Teky5FGkpZX0/gjzXj5Hjm+l5d0NdNIYWZIAZKBOh4V0sps8
I/hYlC76DSBqPs9ZVy0rpcFP0HEaQexUQ6IuiQzAw6E1yN5QCEtCwTdveSQmGSAMOEk+u4drgUpE
o0kYqwYWpsgLgusOQkl//eTsUiUwkfQ+LQgtGC8cd+QZFj52ZqqnhSMp5PP75wYt7oI4NmKKBq2E
I2Yamtj11lvcpTNBjHqBMlEUIUIqPRxWY7PwBrdnd9P+ESQZjDDfX5eomGBvGQy119VAhMRswpgf
jYvrwjky+upGHRtsCqR7dTprpfSujusbyquG82MD4GnZ851PGh5oU1Qe2L9A0P7HsqVK3Ka4WE7k
XyujkiY/9Vm4T241JE/gz/nLqGLUa7z/IbQxj/91UmNP9sfml+3gDJaXbGASBQh2NHU3Q5H+/mFq
GsGqLY04+iFAT9pfhIS2y3hKdft8k61Ufyu3fjwkk6SkKvND4G5qEn3XaIMC7Nytpyb8luDSbB1A
wfcSteGkeURaf5Lf3WlPwjwX8aNNHY67g7pm9ztKqG5rKJoC+0lqReHFgASoohwu6NfRgTlyoNKl
kPqXKsiIZ76ovy5mdyYQGll+Kn5xVZ9dGbcGLFfOUligR85+2lAvKCK23te6suDS3v4jlzRouhTq
u/M8JtQMYNHuM4UqJxpkp62kFcybjdIUytY0VptWyWKJaS1ACMNa5HUxCZounSrZ855bMxm+vBpI
VQL+X4t4bW7SOeII/YjYIOnvf6FqHsnoRStJmIMCeqifaA/3IEvAritBQKN1Rj/ABA32rKzkHAOB
IH+Eb7XK5nDs0xD7yagJ90+bFNu/PA6A4rhfQ/dCWttpth4R5QaD5tydQgxDNEw6Diw1P9qblyWd
ksG+VWU/ba/RC1qs6z0bfkc8c9l9F9zDREZuUnjYhLlR76SHefNuR9Hj3XK4NlEyQ4ohBIh58xL5
vbo47qVTXE4BGT9DDidgvQcvE/z5i1rc2AmMw60lxKP4WmFfKNAOs8r7GrrQ1DmEUaZ26+658oeJ
pdRPBQnyU574CTOZadts/Iva6cz+RaJ3IC+7otydr9edX4mg85qfeEehWY8ytO1BA7+UIVVEvBHv
IYqAhaW3BhAJSTXj90+7OMHvGPUqvAd1uoX2Ghga6CNGkWwnHZ/UFcbtwgoCTXfbnUqjozXb60rE
ixu54yMEu/x1cA8KeuI8A5jvxRuD8iYYanV537uMs0ep/260VhzuButR9DA1ByGwaUJbKpr5bA5v
g7bS86DYEO1RE19nKC/izxEX3b9kAuNfSHbzc33HlmkDnNX6HTxLFSRSqtHlkTiWFzM2mlqlPS+P
jXnFlmkKcZjJK+Z6qgIlbgENZ9v2oa842oF1FYEJqBPmAqm5tzKhsiF13yXNXYUjiU4y4COVW8U/
yUGRn8e3L11UXLXWBzlPg9M2Sz4PuBWZ0UlcV1zuncOAOJJiIGpDlyT8xUZwe0AlWUnE8W5EIq5Y
99BvGxsJ64AzViaEZTa/+h9qXZ6QINJ1crLTeESP0hm3QKp4p6+ByT21pFpPiaHi/OL9VlBXtmUr
bJqh8guXWCOlsYWd/BGqi/r5p8e1GYBeu/E5fxVmffWyOU3d6JlYPS61JxWA9i8IagvtnbXNJCke
od3BfQLm2Rpw9J8sJUzWcQWfvGhkZS5uQ9N6kngk5T62VK6EWdjxLdGy9LFDmkvV2K6fsz9zGaHw
IJE2UTa2+IMAAeCVSHb9DVZn+6MeABC075Ge3S+w1XvXZ01uXt3v+QmcqyoOnXBuobNOQhcmhOvT
BWS0WsRMEw5KN28crKpIdt1Zb0JzklFUCYxrfQA3LyMjL9TFUHtD60Ol588UYVuf/X4UusWviQVY
CeBhQfBGEYyelKW3PfdqiFm0s+sk3DSOa2qfqdx10YAy7W2C8Gi09qFuGAs/VSjRDN8YSeaV9ZQt
zO3t/w/itmYk5iV+/5Z9+PO+veXtb3rNIpXMXEh9XhKRH7FdD/xSh+C7KTRoKGK8Dbv1WRZOTbJt
cJUmscxCK6feLV2tJEoW2pBrAVnfBxbEagiXRb88L3/GHU+hAQy3y034qhR8vvRTS2LZvJXE5Gjv
dI6bLng0rKKYnsguGn3F/ADiXpjqmoDMYH39D1iFt97T0V/Oq/FB6xDNguz8X4W2JF+S4m6AnTsZ
2ZkW8dsJcUAvpUKT10nccmYxH5hyJteACHVM85KvVhLp7h1GXg8QysLabQiyDMEDaSds/FzcV2M9
d2N9y29E4Ql8w8EljzSwNXVcrbP8N+Z+LF9DaCRBekXsrLgR16pYRC04+o9DbG7hYXjy1EwvFWBQ
CYjkOfJ2gZrghRVCiRUc0L+BqO3fsJJjrjJ+aONbCQcR6UtJwHVDQ9jbzVjC5UX+P0nm7ymMykn6
+gI17qdMNnVinuzj3aE4HSY7cndnntFusRRnS6py99GrZbXTqAks+iyVVMGrY1NK9ROaczFptKP8
WYedpqHaai1rZfA9Pkm0unFIhX4D5U+fQLM6vQfkoW6XCIJwgXCtfLroB0v/hwh9uHZZaFjqIHD0
v1XnUNX91pJ21tp659qfg2U+1lF53Rpw8oXt9bOvsLZTPI1a2bwwwQTO/4XWQHSaebNjpUnTP13T
e8wvXqj0dBKEBRivv9/4QwG4h5w9PoX7+zgSAK+87yDGi4qiwc/uIMpY6WgAzuN8fSCyHDAh6p4t
c6jD8aWoA4AE1t79bDWyCXUsXEB+AEHM++J6F5w+S7NbQwab7N2SaeLa1WiJjgF7dxbHgE4B9CPR
kQ4NM5CAwYqB0QVIYXu6wnIuLT1ajb+peJr8MOPLV/W4LW3TGvwRhUReMmCxuzabOAkVT9pj72JO
rv4m0B0IMC1NXo3viUwewAqoY95oRrFdddFF+FrZJLiTV5dm/jF3GMnebY53vjRk8CZtx/ASKYyn
Xg7QPnp+YD3lQlyD52v0Kw8WhpaP4fTtnaJXB+O87M4v4P/3TNs0mBQ4Hy639nO4jtX0b6+M0Rrv
GbZt23tYUX2plkFGyZBg/yyLtURrndTpXcjWZwSgKqOZMOTofZT3Oyb59p9uKyIBGFyL8eDxKlRG
CxucCtsplr06AFL6Z6z6hxn94cWXfAXLbeV/6/vXfvjBLs2tvupmkEVxApuEGHBL0IxK8TcJIftz
VL+xirJI+EeVNdq8bFUWfy1/q4dk2bY5zF75WjmgdF8gIo1D9RcbhzJO/dNGPNf4hWuINWQDgCoe
Q7ny0HNEZ2bqzXz9w+V67ukKWtxpQKJJxniP76c4DT4m4cn9WC9d0F0hdRQaNyp0vmN5GtekprnL
pyXIP1WHbURDt3EbFhCTrZ/xPd6yij1VhJlPP4gcnIpj8tJu3HTef2+K4QZVJrrF5qlDZydvvW+q
jyiiJR0OGqdrVUqNkLtqQmbwtdIAAQr4m3lFHjU7X8k1aH2EAAaZa5NIbm++czEWdaMs9t0+Pq4J
PnoCkaObgeK6fMEDW8GD3XtDpbrPRcXAy+WC0PARzZ5uUpiiJPZZ6y7hBTyAM1qHD+MTK0/Y+Mvv
p3goc0D9E4JlYuQsJ9fNEGgI+fjMzP5i2kMZ3DLTpaIMxwnjzEqbQh7a4tYl2nGfhyJ/HOsUyP/X
2piifp/waIqJ4SYiqxzycH6JEO/NK1GyjkBaLWCqmV54120djDCe6l1arYccKLL5EvW4Sfs0m6fq
OJ5yNjOujM20+OtQmGLEnr9UF26nbAArBsqYtq8hajvrzAXB/HrO4SzXc5wFELiRf+JgVl/0x7tV
/lj8tRuM+gBp2WH7yyf6S5raoT+M7eDKvXfviHdn/oGeGCbLVhMfn7/rRuM44s0yV2AHc+8IYThF
Il0ZuYyWw2uMz+fzTzz+OlXNk/IwtgQauCXd9dYWrjsG0csUNxGqnMxOdHXEOfiMMcl898U9ZYzy
mVolS0U2jY02aQrqQll4K2EDWNbvPEOoFfdTgS7Mf/PCY3ulIKAZ79GwG7wNoBEOASuGSXL9dCFI
MEBAIH2RAmE78437DXfhNLhX/61Aq76ZVtnY9alvHA+tAaDaSMTwwD21DTVFzuKsUKEzwwPcTtsy
wYR0AZNgdx0INtNb/iBFkrfMd62+l+bIVovNOYzC6Jv71PNwdRhoc8v0QIxu4Ejr0hpHbUQn43gY
0wrAkN9euqFWRYeqhqrXkLecb5m+v4KXGfzPxkpG9mTeP5KO/eOfWgiBp7LdMAy8ySAy5uwLYirD
tIBrLuwW/OI01PMoeogEYD8a/8gzT1uVgJAH3A8uOJhkfT9DOj1hxy4L2+hFefbPxMwrDAERqsQz
yTd6rRDcv5VMuIS3HQX/59LsQ1EZ05YweUxRBb1dQn7EUjCjL+KaYXSwbuMEJVV5rpxWvkqhTL3+
5LKoPJhfxBqC0sKA7GgpGyHPqCytqpFDMwcyh3a07n1cPfLvVQFqlXl2uqK8CoFu8IwFsaLwOQym
NE6FHtsdWaYutKQ3Wztrfg5IxjO5DE9nqedcvr5BSeXyufmslFelCQAd8+EhHButriBKCaFzrGHS
tDkDdcjgp5NBXe0qgAmM4lxX2yzzQSaQ1mnsVYdVblLzdiOSymlE4qTSVJPzMFlzWmDklKl3+GW5
7wv9WX1VSnX1zBTDVTDL12iuB6gV8qJGFGSwf6bpvzNJj5qAs7fN0tFUmvln/0wwpud+WPKuQhi2
6F4e8eJYbraboYnAjWdKN5y2Flo7+jKyRx+7nCkqGTEn1gfpBWJaSV7Ezx9xCg3CXTrrTJnyfuSJ
Jn8gBwy+7szlFjlR4KkFEuRRF8PpEKshVJ2TxmsH9/m5rw0NzsBk5jDb1TdiFxl1H1pn4lQojEyc
rpSRUisvNuXP1lu0hvfPHd8yNt3ccp6C4JkqbjcCXmIXjeHjetO18mVzy7QU+YYQw/IDZ81G28Lu
5VnL7sigLykQXjHfh8G05Ys5+iSUp89De4GOs6xW6PDDD/xsnKWl/bwEpi6ahCTIn1zUK0vkfu6R
SnBKHR9BwJDJAoYLSfw/jv6XMTxdHP80ehtWhB0CQa9IFriavg1wMnb1toE2Y6B0WGwBjquV3J4s
TJIBu0Nu6zbnP9wkw0NtUqiCAoAnoD9rGRCeWsu4Jm0Vd5eiwJDpCPrZ8rTmq8ukNeJGredWo+Tv
sEkLyBOGQ6JQYNU34b4T/fjH5utcy0ivegWu52rBrpOCTEGV+MiLHIOoLXl2UqZVZZ//i0Lu51JX
Crpb6dcjCo4KQnvj5g4wzOH4Rhfo2v+r4/v+O6fIYCPgSMAlwWkqhGt0wGBYFsPHRzs9GKR0Rq/3
5tPtFQJG5aGdWHfYW9eMuJttiKgq06HpbGni54p0LPNG4DdDWVzPdtsOpTbZ1TMC0VTiYIiSR9l7
sK7w0bh6yoEKfh7Od+c+tA3iBPwUNT772O1fO6pa6ABZnI2Z/mAdDLrn4N51osxD3d/7//h0jW8a
AWjnsTXTmCprFijerkGS7/rvQQp1O6rTF+ivrbzUO7tEtSFyZBNZ/TqlaTcSA5cCeV1mT+peVFvr
hfZo2v1I0gBkr1P29GJKu3VVzfMQR/2JyUzK4gIg1LBC0+txRoW8WP0Xfatmyc7z7WGz2hOqBJmd
PYMw09uKROD6zOA9HHBm1XWgKEuJxjhwVfnStCc8Jjq6T+UFk/WmGcbIpvCl81wnTX6DUmA0NrQP
BaQXOvxkd4frdBzHdt3LPNpfXjKhUGb5QFk5f3RSOCri/Q9pCNEjX10i7SBGnOSLc3ZNFQom3uIV
4qk9G40z9O4OfSv9PQ2kApUFKs93MZz+h7uHbp++lAussmAOHNG5YfOMMngnzqBV/V/MBzFuM2sU
AKpnQmP44APFRRttKA0Ro92D69Q5jM7iBZaekYLbhB5I6iEav13zAkd4ORojCce/ufvnU7JJpots
ynDIVl9mbqU91V2tprGTM2zp9sfSVWpX1Nm7E4n9li/2SLLfByNy/+xgIJHogRbPqW+Hb0FbITgJ
am0ESH6al5lkRLFLLZwzJOa4i8FNx3VYWS0bxBBdg4fWQuv0hqI7gFBA9nQ8dsJjxPJRIilbOCa3
EnTF9f7xza93yvE0StJ4Me4aXp9GVHzs60RwXyXAXIe6U8kNqCtqrF0WfVIGcTT2Y+X2zP6N7f3R
+kb8TAQrkCPXTBbXN99oixqBbS4zIfs/ClS2TjRPbRW1KUgfXuwA7XVcI8yMq7XxaU4EI113Swn+
l1g43I4AjSo2UcudprWDpH9ZB3CRTQHd7D7rPQGUWJ5PwvslbG/9OyYuoqWN8EXDzPsaN+vK2ghX
vA38DWRdtd3bsncKw39zuHmYtVlDwQWWeyowJWxIba6zQxIPVlv+jnKVD2DWSwAlIOhdQN2w0TO1
n59wDsEnjhPe4VJlnQSnoa6Q73LP7McsHv/KdahyApbBNBO2uJK8B/ELAsK2xjEIbeM+E3J189rs
ecnn2ErJDYpY00UB358wEZCUuw+Mkqpu+A7rnU2VqK8s+/0UWm9YdGoLcnwOdGBii2b63RwFVqh4
6zvc+SWQamWm7NWBwNAIhS3MrY3g4ia1ykrTePzrhlsIpNjayOkwGVIX+HMY+DWXXuBzOPSX5WYs
YzyvyR1GgCwGF/aRf56UR/ijQf6wa9KQ59I2CD7iaqnUAo73q9FyZittfx4+8Y50LlWBxDG0OJDh
SVQ3nNHmvC+xEyuThTafGbR+ymbG4XdmV5g6E2HLxKe+dK4hEpWUbzVgWaKr9UxkGb81OGKWpg6o
yW/glQVgr6kzp1Xt1871EIo75DrnW6RGRac8QECegRekOIgjll+2LZFGbyhhoQhnwSvb4FKqMG5j
DMwg6x6sCnYYq8iGyeov9iXtS/4NW9+/K9UOqPkBg5VhcOkdTNLGQZBmdwo9jdNqkPsF9fFc1AxU
cxSJLrBoMjZH3E6sVE26A/UUajQMVuNobo1mXD028xPOXlOFXn5ab98e6JiZ45VmJwjvrQHtQ3Mt
Cn3EqnOBcEReQqnswpHH8aU9tKQzfToeyy1B/DODlulxK5CjaSpiv1zyBtxuOnLffupj5vwWmXNF
jF9LmlVVOYF9SNkPunvB46VvZzPn/pu90c6GKHNAolsaExDcW1pTwa6pE80Ddj95NOvzpn9VHVO6
HCOFf3ZI2it0Uw6p8Q5BIGf6M09KgHi7R+DjwGc20GIKT7Y7oU9h+thuLCFVYjcYAd0Mkgr/ppHY
VIqzyBzvhagcHdSswxJ0RZDHdcKefdWuFXiurMmq4lVhGqCuTe3xUv43scZ7y5epOtEOVOudm2wA
yycY37zc96SvqE9O9gFa+MtCMx8L/H710PIbudwUL0+QHrJvjPUCTbnaKuwTbTAl6Zr66ykDNFA0
lFeAmcHwSgqtdbHjufA/AjMI8duTJp8NikOheRspf9+0HVDFCrhY/xbyzZJybu01/xlH2AwzB3Ey
9yzY8qpkA+EED3RgmRPqVcn52yhWi1FYU1KTwFsKYWvnb7WPgrVo+VcNvigPJTFN42f3PoMbKU+f
A7sL1FMTBOXEVOVN4dSw1ESV/AkiVOF++sj+VzXQIAXeK6AE9YFRPfO5z83t/Z6iczrtNlbeVbHm
1OtJ7UfJnNPJrq9JpQOFkkGKWxA14tPnoZvyNIZBCEKaHCVGu9hTT8Pq0fPR9bDOrvdy+MZhE2c+
hdHm4GYmbUHylTcvuzdQd0M81g34PA/DUQWwIDWX8k+bJfTstfBI9xW26/JyG02uU04Xi0iDElwW
7BhX/qtkHMwt5tFa+HXMq4BW/6Y45JvwOkiBCgJqIYO7b0cioFInMlw8zCIwceWtUMJFgGgQv2+a
L3rw5EkKUzl/J5omRglRYFJYSLvdY3U5nUgA3stRehpw+jLTp0b4QmhgdMISuxdM6ofxWkEtUaM1
SpGcCxXS3Lz2JLmoroymzlZ3iRmZPvhHhqYNxD3asmYujFa86SOoo2Pls9M6ipLt9UkRD/wSWvGZ
y7fqTHFZ9oBFNxQY6QGWF4uxSDyHv3hS3yXd9fidsEmWJng2uVdFZ4hqru3h6jaW0FUWrmZHzxRt
MlkiCjFAn0txz541jNSNbN/TEWSPFvku+Bc4R+h1iPwLDE1E5W1qm1nm1a2Bbj9scWK6eyx1CuhT
f15Sk3N7uAmxNkH+dQwmlEexcu3aJFKNbFo6bScECOYTpJRF2NOoCyIp0n2IhEs6D4fG5H1XGPTF
ryVu9mIGUUDtrYEnztq9EBaOjRqG5SRJVO0YrwxQe3ruEnAreSRJwiU3f/KJdZef7pYwdUVpXen6
7D7LyoWWUn6xs6+VpLQ+BUJndFkU3P6zNx9tu5nB3D2QBAh+3KYvJIZrF5mNGsnRRjEmBvxyL8HM
rc85BWS9qo53wjjfOulQFEbWCH+KzOI7KCm9iMb3Oq5AWzWw6UKysNj+agQndKSmubTShXWGihqA
6r14bDWTdDr7qCx4LGbM1kbrvMsoW8UNcHmka1FXwyo4tIQdcENztvABNoMNzxL3J6MhDrBsDGg0
un9jN3WMddCW756lRECrnOuGRwtnlkgNZt0YkFxzGZQ5vUrPe91Qnk7FB70OM6OmxeNpC8+WfH/E
MSxHH6+yq8kdbciADgJLRBZvUuPz1R/sBdHXajoRlvXDAFvguDWVitH8mBhCa6WwhWF3iGYYrz08
bM0X06txgjisNDA841vbbrcn/5ZCnqTuN89FlrgEAKvyBbMwueuWrPDavcxQHg9YcErgzYHgVpe4
hcQPgvShX0gEBxJU19T6refA1gvWj7QS+/U8dTk7YViCVC5pSWjVNQRBcJ8Z5IfDr8vfCgwB/35n
VB3UfYcQarNPEbHKTo0LGj9/uZqqkRe6F81NIEV3jUmKd48jJi5DWgnYF4wDRNPBaGNlidqQ0hj8
wlgvjhLjoxB5VPGkNpnsCRN2xvJO+lb6jDLDSrna8zsGUcTvbWvdEbsJuv5Lf199W5ccJcE9mOlv
M4X14h1vdfG6HQ4H3HYLvud0C8fnNjEDq2TRLaKD9MbHkV+aLeE0rnB4D/ba2GBo4NVIpWILtfBl
fYzSLUNuI5kQU/h3+3SWOzOJY/91JpmwvvGOkKK7nGx8GtpEvMEz/4yvbqCnoonA8obdbZKY5R+s
OcuSBjERPO7VPHiYoIpVaNMJBJ3jYIY1QeobFcMeGG+aXemgeuDLFvukCuyOA7XSXclizNMipiqK
MU1Q9rzb9bqASqJgKykaP/gb/3p9dzsK53XbugEQoqhQ2gwjyJ2883aNjyn/NvtokEUkzwczcegb
SbuGXJxI+6R/+2vometTKXZVBFx5IoVVXmx9SEXidLV64e9Ozij3EfxzWmNIas8R2EetAwj9E6la
gpNxhE3dv2GraXQhsKFstqnpcMbDV+MUqSjvuXwLRHZyiCMw3YIxyUhk2MEjAIU13BmnSX0qRTM7
QOXWfhcTT6d7P7tq8g/2eM3jwn3FKo3+62h3Zt+FjQQ6viLvCqH6H1jT9Zmt8P/LCPGF2iPG4Nku
GRppGMXAh4OmLETxQCRN8DDgOoaKWxx+o1Zz8rDRmK+497BV/kVT5C82BNt1zPFJ8BKigvJY8M6H
DsXNp+Zl1/3LR2tIBTFWmV5tjInQqlRhMTBapygJTP2KOsh3p0TpS8od47W3RBeIvO6VeQAiA6CZ
WizGzNbOtBGCxD6UCxny+AdQTBOhuT7emqBF/pIw1RvC8H3MfUajooKYzKbdo50V2uEK0FG2A4D/
LbOixwOtnZcuqRDAN9MPArGEmjnVILXAtM/FTwMXdKlys6EDlk8UBBKhl3SCbNNTjRQdRPu7H0PR
0dqhxUNef6mHC5c8jVAzlV8q2D9fh7Lenc21E11zAiwZd6tXXXKKO4wzhDsqZhYdK1saLBDW/xfN
ush/NFmRm+cXl+uJLUOX0Dh7nsCjN5s5CcTom1f8bD8/lGqmkJiJalJaTKQe/jGdKeKOedpiccfH
jLNaePRud723UVJNAUkRQN4SkzGpGuSDj32UEsszPUNyi9ttxXgVqQELIKN1MS6YFkC+l3ORyWqR
uKVHHoqX2R525p6Gs3xI/zAVLbwF372rWZqkG53hYpetm1J9ISj7NvkrVWv1DjdLeIrJwNFEsfwa
BgmciLASBWCsbRkezX1p8hIjEjJZK+LaIduOne1lklWExGHHuqfrdV7t8ex2f+BAzFL2nQr6AMAe
AKYp6B9nSP9XVJ8b6S3mKJYbNxkYotXHTtzvDuvJPS/pemXYo+sG+I2JUs8KPl2uF0hwi/YK5trB
/1Gu/SxWpuzxBNrNeWJ6QiWyprf6Jz/PopmydK7gED/GWBci+5xjwqZnQ34EUhehvDW2fnWE977/
4gk7AdcVSWIscv0t5dEYD5DpYingMqW5PxOSUYlAc3tuzp5sgGET6ODSovai5VBjsFOF7KERDl5L
i9dex7yhuObA2W/+6ItDw6VbbzzOuRdVA/638x08t08xn3mepsepmnahmS82gN8pi25gUhtZ6Bw7
miGk2rFRoe/bVbR5ktwU298jAR1DCfcpTqDghrP82EDO3obe1eGhu3WvCCnVymTH6h/9EsoXW7VB
IPFjUnoB8ieXjT0eedpnUzqcI1KTOfAk0YyYYxFFt7InQ01i5kiMKA/kjO4l/T6PXZ5iH8UjLOg2
MMgqJeJsZDPu7jBqpkzsecnRhchfcGBeIRpbsG1ju1MG7S5KKKXMT8uHoooFNBRWo0HvAdAmW7tN
871aIBLCAs77jWdAzlDPvpi4V/2xsu5N+i4ORtbnn8Y0Lez5SxOVYOZ2pykev6MBDqEFKVsYq/Az
OnG3MUffNILUb5vb2Qr9t+y6E/8XnPALPRMFOP+weGx0MTOcj1Pldc7zZ3M48n1SO+HOTk6DBKQE
BPiMh+9c2LHR4THZFye0JIQtZZtzIzjcH1fkVzO/FxwoU4kyL0+rIf7t4nYlZpqWDR4oZQcShC8e
azqkmRXEJ/Mphs2aguDq+fq892hlE6Uy80yeBoxx1UmkvVtGWzq8s2aBeuoJIDTOCmcU1TKT8y64
GbzrEr6Rz45eq2SbvIclXX4mfDunVAtMEvVrNWaShmwzFnyRdoo1KCzFtrotdVL2bAdIUw29z4a6
ONJwlveBHSHQT+oqzUqAx0LDyMQ2kVQJruA7i9bRSgBD6EbSx0ZB6AOKwgWOgVOvCS5KuJbdx2/U
Iy3+Q/wN5wlvZ1rXTEyCtkUJOTlNyhX7nNG4s1LmVOCjPebgzMpxVQiFZrUhAiZ6DT8LOvBHYe3T
F64SBDg50T0nLHwoG1cDAHBT5TKi4TwKfnF5uV3dTOl2y1gK3rQnUcnUY/mSBBhL3CHa/x1Nq7+6
rOL+xQ3lHPioPVQI1/9/qrWeSXatU056Pgt6IkptZ1Ks5i2t51yxc7u6o4JdiPCakEPtVdZYrSqx
JDdNeTjsvVt1fhavsmJNKiwqolSHPbsa5tU5UpGTAth+07V9mnsAiEFG38KsRaF78zpPrpFCnz6r
5PSVI2mbcw3cSt99kWI4RZumqKWBwhrwhqAh9gtdADy65xUYAgmwSBwSAHtvqWtpsXntDk7jP1fq
QYietWCicPLvCFWPnyyTytR3Zoi6l2e8PnsCi8I/X8MEjd9IyzuCTLfnvXz4LDoTmUE5q1jDrHFN
QC6+4a9Rxx4+/qWlSTu53QCXidwLWvC5RiSM56VjIxpgifQ/9jEHuCbPw+l2dkUunvmSNSsQyOx0
+7QoLf41339LbgwFjhHG1gV0Cmu3k/GMihtFJHFIDbyTNPSbZajmyparWOHlAAi6r3KthwK8Wj1g
592Pt1r9aLWelN3qq0UBBQ6gdCaLbKPabp6TtqA7irrE7AeiscAtwkUVbJKZxGANQ2LEe8p+p3oC
uqWSljScezjic2GE6ZP5bWo0gKT94rZ49LrjqqUr242GyPIb0XaxPzkq3bJF3xjRxKP2x/E/JX4y
5zMuWyP2k4shmrISxHL2ajOrWPtWeBXDWIGPicZxseHTGygM54pdWGBSoz8zs4VlN5cwJ84osGmR
t+9tQWX715Mi4ZYgTn3XbEZ09MYkhCGz0UvmfPUkR0T970V2muxSPFPiIemdnqqCrvv+PzF0Cx46
MHgcmfaDtYIiEqRmE5yzV71JLIwMkI+j+54PxYz0l17/Nnhn6/RbaB0/FgL09rNnu+mRNYVI9xKo
Rh320RrFj1gdn04TUTb2D01aQ8xoyTFhLQ3Ah+Yk4Xj6pqHT6bCMfw8s0G3H4ej2NHagcyxKbhJ2
tHZxagK+RMWS8/KKvEHEBviQdW4Jhs4p+6R7d4h9lqDb4zbG/DSzjYeLxM1sSWPfDl8rqSBom1Il
tID6AY2tD8XVXFvDA11xZMRH9iw00XK8FIIjTXQeHyQXMtbgf2RW4Wgr/eYvdyG4fiiGtQrDhNXn
rxM0rfGSHpYFTX/fF8qCgUTexADExfphIXYgNgVZ9MyqjYek4IKFFgpWDhZKwIyoMZ07Y4eCxDgo
RbCapksG7Rm8dihNkd+vO4IvjMpb3U2W2BKQHMXTgg9KrZ8v4uYk7VAnFwF532UqRwzY2NgNQUvg
f1u5/f89n1e5FxkhgkDIwlfKrYg6d43IPa2aB6m4kVCt2XimTp0aot/pSmPv0J4UKd1Cwxr8tuTC
lAKVY8bSVZ2ZyD7a+ME6aYiCijNR/GYxIHXUlXacKg3TrW+CuOJpGk/QyCKVltg718+6g9eNcSlF
ExWsMFebre1keL3sn4v0dNSGrRIsytIdtWrQCf490e9jo4o5sojVY4EoWvZXbwzm1rNqw01FpyV9
bfIrWwpGPNl+qfZ1+KWikhgCDwff/g2LwJy4w2KF0mAx8F/hM8CQpct9H9O4thKlXQJbxl0+X/zg
Q9UwzsPVJEg4XiE3pIZ8Ivpezm3LXBN3RrW7Dt9qbDDnY9tkn+GvITh1NeNX6mzBDMcDlOxTXS7x
yKIoaarqjcVj6pMP4bEe8BYwJ/PnwT5eYIqkBFOa6rj6KQ+vAemMfgPG33+q6lI99NknYzk3IP3R
Bo3h18UUILcHKPo2vZ50AgjelDiUFZK22gYH8005ALYkgRXE1HBv44wTCzivU5D0cNCPIjAxGBgD
rSRDv2WqOgnO0jbsaoAilh9iQUv2HfYISU2YjCgfr/IQ3LYyVlT8WMVFxkb3ixQzGO+/blYeTH0u
WzK/XaeZlOL2579sCREeMB8Iu8YmEJRQdydvwIdHTDFaDcy6RhzVXdJDvVETpx7pA+pwBOkq3SQJ
2Le2ivWUW3y3oigr7Gdp0Vvnx7b2godyw1GvEiqsJG8Sn6eh7siRAjhmslb7jUo3P6O1Ypq7R9tu
uzDqaChYArwDapKsfV9kxDEj1Ht7pMnB1Hl14psfNppJbCxVg+isnaVfh/Ei7sVCwU45vBwnrFdr
9X0bjzk9lDtRZJQrj5nt25gQeheC2EOn59zzMW7M9wNnalMN7DieUgH642mxOxAcQ8TiePbpj+5O
gK5W3ChvizEtDFqKjJXcF3dDnYmpsIXCi4NvdOLFADBvys/7y9GK5ebIne+kkmPDETQQVDI1cH6T
tqpx3v0iusCpNWLXFdIfPbqFhGbEwmaIwPoM6zthMqmXOfhggqKZfhy9KxvzXax+qIJaoBIvG1L3
2Ih7FLqlu7CJeHUnQBW413FvyTKQSdDmr4x5Ja3R4hyx+ReaiUPzazR/0N+oUmkANUezxMHRwXaG
aBsT431e2vlVuEf+ANu6nyAvOTHtP3Cw91KWetPW7ZOxeOoY7VCSI1pdYnbwRVr/FcXtl5IAxJ4v
cdocvXfE4DMjU9quRcd0aJaKWoA0nq5K8hPKBZ5E2cSO+eG9+iBDXJWy4ZwgWtwbBV5luK0HQzMB
4dkoluAPKxHePGI73e+vvpPSTlUSPligdgdqpHeLfLocL0DppOUS450EzunTE20a84GEQP0duuh+
Mef4UJUE6ITzVj2Z6b4BeZdlxl9yaVzyhfT36V7b1tmFnzb41I5syzCWw2iXlFD1gYpynKZOsLEr
ingrjOa5SfRX/vDNSWEN2P9IfSG4+G1zFSSDOoTndpeKpfEkIISDqYpObbFzgoFmri6RhXDyUpbN
bhApqyl3Irq1xWGzDm/jj542/eVQkD/AeIoifyc0jVnHcAm+ZebiPeHbrgG85Sd+AKBZuxX6fxlT
gToW84R7uUEXI9VDIrqb3fRbhI74VJLfsyHQdzStKdItAqMpFgAe4Iin+HT0VJTYjdOBarcPb6iT
HUwJHTOUBrAuIhZodD2l/ehT5XPcQ7+YYDzTGHxyKYrLbuxfjjbPRqOKTfIUxmSHARejBJfIlWCJ
Dr2yZYy0TA02pMVihdAAKJJVsq40V5XHQlCZ7pXCs/oOz06caak5uYzAJsUqa//0HmwK29Le+Ym1
GSSWGcVBY4xVnaZG8j23zJFpRd4+iw5xbIS3Io6cKIrm1fS8U0c8bGVJ0CpoY2zkPwo+QKQ5LKpG
UckL+ZyVaSFQbuvpA9BEdc+VtrBBMR2XV0ruHo9T/pKc8xkdSx0oUrRGM4gIaqRXhFA9n24VA2N4
frBXtcGUC41P7nxMz4eSv0iqMoaYgt/rTdIcNdd8D9w0XiJS+xPbwMKMXdAaoDvszYwn7Bnjyh9b
ZQnGCglcysF7VxmakDBHIAA1F9kx67twKJC1uKCff6Jz/0xSSxQlf/QESpsAIyJLzFs2HzA3j+Ny
TaZM40tt8S/fPd0cuiUG6zcs75VVpVw2zAIp6lirAATDa17lFl+EpomCFQiT3Vvkryp7wUoEIbSn
oe2xofBmfXJtq8JK8w0/Fr1upXp6wHYQPUTZqkyjlkzC9zHPBVJVC8w7pKzV13VX2o1wjZaf8Ffy
BFW5S/Byg0rNF1UDryHv6owNCw6nxVfW3uCnkxa1ao/WqhMAjrk5/BjWmWY1vX7QEyAI5FVEFwwQ
KuLi4a47yXPtQBQ4ScUBKob8EqEQUz60vS8aNhaspwQcvHVahyyOYhmXQW9M0DwYgaKQgaEX+E5d
mDmWapg1LvHhfUs3ultrMQWWDjBgh08MTpz7s4RfduF0pzWqN5k4GaVJ+pTtBJksgNbvVnm5JVP0
CfAiyW6ewXXuVYH8Y57xTa76kyuCohdW0D1krpnuciZJj10xcQET2/yk/mTUxOOL/xldLhDmexSS
Cori3Y1cdU94dCnzt/gQyPjwlpdlBScy02ZFv8a4FR2AS4NeGbX5J7DGlJcACWDCCmjCdiQVk7Ka
WC7tt2bBpVVE/VwdDEroxuDXrd/Ne7QCm1FiG4JghJWCDwqalkVzhLXAHnxcThcQTVhKw4o6l3hs
0BH6i+J4t0a+KMUIw+4JjoCWNAd4meJCoSjhvcrTOXWrFprbObAn3lrfHvqz4m5yNUNspxlPMiuO
c9qsAlZIsYZU5Bcl0bLkOCGakd8MQ+FBnjtTFCp0PACE6cudjuWht20plHbZhk050k9gsGI9L3ZI
WEHAaAPjZONX8lWbxjPIDoAsXbVPZtb1V+mWGxFWR9s8fRhfeCfCphlIBLZho5NNj+4AK1Wf1fTu
0/lUy4KcP8b4C48cuaZ6RPILMcFypo4zSnqMHWz3u0LHk3nFkfwXx5pzYXTXvji1cdRlpfDbyV2Z
Aq1M9FxVlkLzZi+SYgq8jCduLVJirV1BlhaRnfuUI7k7fIX+8aMSe/VKcngS2fuMydHEOFS1F7xJ
uzcaXluqhFY9dN8WNJZ3oR3t7LuvoacxgKROtKfO3bPlzDZbwKUg1GRJBsV0tLO9Z6PistoKrnaZ
kSLC71v0HNphttuqLSTqa23covw4rcWzR/EKcYUFat9U7745Kqx7Rt0QTUxlQd8CrB3vBA3nMGK1
zpXikg0bILcaEqCuCxe7vK8py//HYwtAbxqFKM6sdRnG9Xpbl1VoAJY1vooALsvolu9Iu8P2M9Td
sjeVw8TGas18/SpJXhNUE366z6hCLKBcL6JiVi77sAa4nKnh116wtF+yf4kchOO5gLNzcAkQ2fBt
SVudS5zCMX9qJ0JFR0+PzmVP913vIQbPrdV6wkr4Vqf8qcVjAOs+tJ7Izl9kqQTMC3t3qEOkjilu
XOdjCTOa8cWLTx1G/P0eyDfVfKddKn3r2TlTG2tXrVR/hfTmWexSIm9F6Clnq05BSrqZ9azMZkYL
vw5aronlnAZ/yiKnaP7xPgD8dR5OxTsNVWTEn+XiebbJQIRRAOwDyIQvWEYl3XdB+z3EejwHAcnZ
fghiJhEEjN9TRjkcIrEIf92fAMOnj4oFc9fW/1iy6qLCDrbY3wvIj9jzerteHEQO/P/Jh8mstDr0
1ZOG2OorbFfNngfwNViLnKu6G/guhIVvFkHiugALZ+WXPYeHadk5LUA+MBTESehUxivYITO6qorF
ymJrhTOU3mzLDIv27xRWSbuKm2RDCtxFyCPCq7Dzhx6Tt/yLSfj/zB1OUQg0CBIA7AcOOPuC0PEJ
Vd/ivqhhCZZ9fc/OcEOwuUVa6z5XAircU6XZrL+fb0j/wEKgCyn4uXm2RjzbSGdqZebtR7ceuX34
Mtn7U3Bqlzs5eXhlypyKivdlUEtQGHz5Sk22my0ZSXRySOWK5bTz0sasLmGhIiyNJSR3rbPwp/mQ
Qmll8cBBoVZevuikxi/ByjmT9ioN0N6uPWNih6+DQWfoEGSkfyEeFSssx7hsfiy0jexrQLWet/Ji
EkOZtZPa49lsZynGHeEyWy+CvdRKiB7qyfV0BfFbFsRSK/x1EiSexl0naWlYmDcKwvHdmv+XjpaA
HUJoQ1xhv8qpG4n66/eMZMRU+zdFv+Ivew2Q8BtVjp/ivgP4JzV03GhKYXpevrxCV8YYEbaG/Kya
5ZaFuRfF3SQbQBURdJ++iw0tPKBvG3rkhPcVJ5oKOKeC1lm6IJKM956/Xf9f0fL1Uf1/P7dkBzDO
MqXxgfcMZXx3BGWRfLiSEUAe+Hdc23j9jhJMES35TpYyayH0wiAkGMjSf9FxLNi5fbpQ+y6V6+6r
2O1rS14TRXa7keYVl0BHxPEP9a/QpA8bE6gvM7g2Z8BZk2WAitPOh7800/5pUgvPrxN+jiIQ2eGG
PE3uPoysVW0vpCRuMCdYKIDFEbJaEL+end7celwWoZZAsRZylma5SU0QFoIHbLoJSQxRX69XHcxe
vvgRV7550/8SeXtHAYn+0+/B3PpEGnv+LvHozRkcGiRk0d+ZFURi7SVcCrZMnHIz+KCmIl8L44iT
8yXOheCxIYnfQZGz/IiRPfEOY9/O06D6ldEy+AILUzvEGjub6BNvsWXlbOfvJlj01BW6WRu1PoRs
Bxsux9FHFFfs2WeRflqhLB4WRVZi68RI75FG9BaEd9YML2PY9F5EXgWdtFxnOUiKJdy0NVMmdHe0
1/LlF8QeUIrl0aCq6Ut46q+Fad2nIBEbFZ8LflZYcfc8dj4QTgd964DMEErUSnx1tYPfdHB6cG4X
cMxRI7UdJZEgo54FmIMdPaoHN+tG/VqXbzLdbOkXgtI/X9FpUm+mf2hlTSjhQKzsreyAl+X8rZYY
Jmf4qgN+YbYAzI32nVEX9o54ACt+h17H1YfhGTbtBA9xKee3CF6aMExLsy5OMKCx7jQbXR3oQtKq
YW/pn8VogYRH4fTY8Q62uQvtgNpBa6hdPna1dUbVOu0GWeEgL0lf81ChL2SVaFveRCrKoWtPaRTC
WuWdsUdE9mUxieFAaa8KBscYU12Gy77sHp6t+6D76Wp6Sl0Y01nTZk98Wc48SBQgSPjdhr+zxKdY
NO9a72bSeqIwZw48Vvo51o8+kx60y3zssPjMnCYVg+oD/fns8SFmuP1UnhaFUP2PxJYnlXLdzz1z
LhQ/pQ5z3zWjAtBv4+TlvAJX0L7DjugDxPglhEPkKAJLIMosd77Fw0KY8K3gY1FsUN26wLXE14Aa
uHzk2X2kJpQG38zIIO0bxRPSZtHXUstZvkHzeakP3NvivFHWPFuwWQ7eCpAtd67zPWdVnOF+Ubnf
464ZM5dbWEbqXf3aivpy1nGB11E8wSjPgnWOuAZ5pae3b5w8F7mcvGRDd64IqnzneBhSetOkssrZ
BOYnyIFTogxk4PNqegl08JPa2C4ZzRaacsgU9FHT9tupzuz1rP3wa/kTvMvek3juObP9rVmTvmGv
ucWknaDw/OWusP9jhTRxhYdZQ+Kw8nyzFoyar70/ttXPK3IxWlJwP2vPcXwEe1+h6If3wMmbWuIY
sH39jbMzYEgxJvEAHWi/6VzF9lbsq+NK00ahlviCaKWSiJdUn39wBenpXNn5b6aHTDS714OdovPC
DLtO48aVPAQopdr/j06fB+rcE4Ge9uzE9W85E5qM+eqWe5grN+NuI1JMZWfqcivewhmYqKsUY61x
+0A33nbUbdsaUIAXeSBqTHJMSSQN1wrx01ZHrkVvmhZLJNd67RSOI/8/C1hYsLnFifXjPIRYHAfI
w8Tu/cQuFXjgx48LrQ21k0kK4DeKsXT6ioT4ETt9dVZ+oeOfuWal3wyW0pVf1KPPWoFLu3c5ngLu
Jq/wa5jcVmutF7AzVA2yyY2wnzRjNuuvxOQ29uNkEELcK/g7mS43dRjppKIUBtt39Op/N4mdCeum
RAQs9YVuDLTzdqeI+xzClphxSM22WFBpwTJBKDTLsG12yX7Re/Dk+rccng+NDK+l9DYQnoqkqcqu
axqaTxGqolpEbcpzuD1w+gaGPgjrHC4MMSPjt/E/IV7NUawCV6esz8zfY67u+kX09/HtoyTdDvgM
MEx1bWQuEAkzpPJC04a2JYeWdwDO3+066GE9ALrvmwLNvxIUkZHeRy7MpCtw1U9ihO8PLglsEAFM
SZ4WvCbxZdR418oYfoSbGi9i33uBtBaiOEHAckcihLHq4PA74riN6GCh7z7yPYQvs1PDyVgZ17Yc
eGtAHE6Vg3WG1DC/yFLf6ceMzc9FSx62/JQ9wBtfmADN6QsGLabBveeWLNAMqrBhQndIIGl3Icsq
1qF7eSnGNMeiw9Onp2pVkoFHubKbcSNfzhkOoT7g3IURGmyvor/7U+K2IpaA+VWaBrl4cIqV/qGg
hpehwdkdLpPYSTwiGwHSmYSNmMcMHrLjr7YTYm4ooy7+aEV0uXzLrkejhP7/HOZReZPb12JgBLPl
RxqHm0n8v8VhyNhhYZ2bRMqXKqazsagWbHRGmFcw0sCmUnHE14vTk3M57FT3QNE+EH26zpTnbipN
ufYOaTNmcHU4/V0ETJR9PD8ox9S6Yb3wsATnm2Dk9+TExoR+2t0iZ54Tr6PkKQxjNWoigQC9uPoz
c9VC02bakEfQBaqZHHvzs1Y9HbXuJza//RX0VjALEv4TQ8PPp/3xM/9P7IhmAWpJ4+vcOj5illrS
RV8Q1owvntkd3n5sKB93b2h7jSMDkkDvcJYDyzZGliH1Bb/zXwQdpA7kfsS1xodAfX50gEYc03Nw
Z37ypz506Ky5erYT+u56UpA7LlPWehG1BNB6inwkW67Pon8addhVyuMO7AUCiiYKU7+LIpwaD7qy
ibdHKhQV6Rs5H9u6V9bvXTa+GdiylUfht/Hg4yhBdTKLBtzAND9Tq0HzosYGg31Pz6NtJ22+RffO
ACuhehDjP5W9qaI9+DOE3kdKPfiFdDYE4xLf98N4S0MymIkWHw+TFJw0I8z73gT+KPeQt9vgSjQQ
1SqiMgVqu0g12T8nnTD/B2FSTODLVcbbqRTCPu/PjmqdWtwZCBBW7JfIL61R7F9zo57pzRMLQK48
Rn8IjDoKawvJB2FOt30jTOhZ8vUTo134gJG5P6GpiDKbGcAI4saanGcqh5lamyCypIM/QWjHVgWw
Un2kTyxS+EiKFAllic3D2DYuOMyWHuIKivKkbQTViEl3XN5X0u+yvLhc6rJLJT/0uH3RJifDoQxh
V5rTAjBL/4h5tc7x0lBgzURcHLnB3GRpGCQ62lfjoxQQREnc6JmZH1VGRaYLrSNmhXv4z6Roa6lL
GFtCEW8SEHEZUBk8aST+otJy46A5eM3BwkitdufACEh/j9JXJiIv9it08Js9HFwp2To12PsZjJ42
6ZbpIxD/hcmbExNNW5jvSVLQBkT665+OajgSHel0IKX7qS9NRJC7ZJnmtk6JZuvvmR7YcARu6Qw3
2+ZwiobzzB8pNcZciBpl+VA7e87CqqTGBMUKiaHZrmqFfmM8YM3xjBuWKlanoY6wHYLRn4nnHfwo
lxDU9N48fTTMKrXzj59TLUFyMDMKd4JN5dkYafAlUEeGz95fbWzZYGB7OFtkdHeKGTGIP61VngEz
u/x43SfKvUFKZYLmG7QBsC2dzz2zv4tDWAB6kxmYatROyB8CyGTZVfgwHljZ+I3srnoocQqmeUoQ
c5roo+lOfFV1eNkpL4oML6CyxoVIH+TKus0LZNGOY7ZAzmjEKmRbQLpreLAp5Ok8o8P1MvB903kB
3UICIZY4bp+9qgJiMB3F7TwPqza1pU7CBVytC1f8nRn+59BDxtS2PzpCRD2eTHPerjr1UXBb+N4u
jEWQMWx8cdf+Jq4tMmIfwANTJcKc5oqKd1XF8csyDGRyY7w8wuFGRmPNlfDm0laj0mNn1X1fq2gC
nkT9JFbWcBi8hlkLVzWfQw1fWxy7b/+BkoxZ24r459JPK+nfsmtt9YULph+Tf7LO4qnA88CtLHHF
oyue1JhNmIsjTwcw48keckOTsAns5BUzH22QSwV6WyjssWlWV9Tg8cICuOvJ3DufN6q8xixIogk2
W4TzWY8ve/UMMjWp6jglvr2R1Q7ieEvrewdo7Utq19U9x9o2FnY9R2+ec6r+hKVHDSsXv5unEX5/
uvgtXRIdzjfaDFO83OHAVFTJDgVRsBUtzLxvh81Gayfr11wJvcIOqd5vwYeLQE23+BZafrxL2ZwA
OVU34CBIcT6LjZygW59EVHBlYH/S7FA133hK+bNJ6CLIlNTTjrH7ziZJrtOCD2pyyCHf9DyXM0lw
x9b0JtNKB7+MWQogiq5Ytqr0lFJAiqb+8QZtx33cGrpHqNGAaIIONo31kZDXeKvVultxncZLR0bG
/UMOwigueeOxb9mDqKRXC6LZY6D9WFzspmfX//3K5fyYqhXA5zTyZXWM+4+OmD9HYmosijVc4Rr7
nHNLd5ZpCiQVNyrX0KpVk9N1mAdxHCXZJ+MOsT2FGQBFCbgKfhps7My3UoKkBHOwooLUng8pbz3e
QOfWSu5yiNQls8ZSYx8C5ONlqNUzJe8JnJbVD3bM8eZWf+sqFvfl0TNpAGzTRODWU+L6bjFnY26+
sho5e0X4kq4cBdUaifZZNvQMJJ4uUM6XFsnA0vs48CA2TEvGZracuJcoR27Koc+Orh4ypu7zFgw+
MyScVsHnjSvrwUBfUlaaOcbrfzZPI+eLsk/4CtVgmlWybK3h4/sIOWGNu2Q4YQHcTYhSr2+p3Zkc
St4QU+xWQItJn77EIiBCe4rQriLHc4KU1OwDu6nAVQ1zTM9PLVmJs/7J9ZaXkEdfYy89OBBKaJgO
DEm4vMiJoXLGguSMXdQH26a9qrOAQwR6iEso1pfu8pJZDKLNA90g1slwTofA5ZkYF0wKUZBv+iAA
VpDCGRualtVOWdeNh7TYpX39VLvfTYi4YXqZPHwoXXtP120anKw3VMU/yGP1K2E5HHoFyvAwpkIW
8h/Wk0fGP1/JAYiXj8liRncd3FNlJV5Mw8wKdjlLrDFDhH24MaDLL5LOuCeaD9zoA3S5uw3gEt20
L8wubl6HHHQYe2ZADc2utCHRsVdnby6aiIL2hKiooc3dg8EG/M6WhJGwT5dzCHwRxMIN3E2nzmzb
QrtHv03hhdf5lgw2En7683m34y7BxbOQnu3LGmRzwmLgMm0nlRrIXCVV26vInKVGivEtj+0Syg/E
KAWvFjwCDB/A+VWJvydTNTCHE/gzC+VovNOZJQ64vv6jtQHD3qjXuKmBDru82I0Of8jMou0eQIA8
uFWuQqQOJAYEGNN/+FlEHKrnVbBbzLSQXGIXCc1b2jyAFsWTslHmj0olvp+mFQJlxILFUxPNh9uJ
7yUWsctZUiweeGh0no+QP4y9a/5oqqmovVUbm4yEPtYXzs8CiiiWmYQRTnaTZRJRnewxoDWBeBbz
fqef8LEH+RGgCVKU+99RVL/UNtW7g/iMebms7bUgF/wqgdULEH4FxT+D+h6UX4mIku2VAeDrVYMx
PkYg81lv3um8KSYyBv9ZccjLA7Y7PE5g+lRpiF7zGOtMi97MZFewElUVYwO0JesNxw2TOYPahvlo
tyGDs2oteGyORojgkCtjrAxe7bEJZ/hE0tEFCXOkz+w5DCqvxW5BJ6i5UyMLC2fzq5F7P0lm2XWj
Q3l/ku1sXLe6gZwIKUbEi9ph/JJHwzZePTv0yYhhqULljqER1DSlAQvVIjwHjduLFjZuAl7mMZk8
t8s2J8riwMJkGEA8+GCkZfskzjZouNmy9LHM+GI7tNFWX1izNunQygOoIlLokIcx742Y2XA9BUXs
BqijSCNgt9pyvTyBJAD9/tC3dwHR7dYmjT2j0cuA9B+dr+VRY2GP+F8hAsBB32bN01FzVZeXM6V4
xucPn8LK+EbWuujDPMXaQBfk2AxjMmenyl2UAQwMF7hpGTxbVnM0iPiuaQDTbxvX0qKlfbhA8bgU
OEB9YLooR3XA2f6LdP/6fCqE3ZfyYB1BHLkK21DLRys5PM4rvNvtTCEbN3mq56nCP69w9oVSZkad
WN35VIAMQCC4wX8n+bXqhGl0akUC+XkY1TIoCIzJatH7gnaM/H9AmebEQT/TZSs2hwB2wNbViZ5Y
vCcSA2rvGogOdAMLDe8j/AG66NzuL5LMy622LL0W++5MHCbcXNFdkLnRBb+bE9VazVzGLei+ZIOj
RTD3NKDvkYGtn+v32KsdYlso/Y1Ix+cS9HgZRifhkgf/db0ffi6e7bS73ADwKepBAUoxUQp1Hme/
zALae+p6iV4jZDQcZxLZ09sLo9BSHbB3KQMr/gvsoZ2OnsHwcilHOmpWl3etKTj3D/V+YEf+9XNO
6BONyF+EOatbNcCy6QJzVViPJh8GRr0yYO+1caWA25xAMmYYA/nOHoCbg7DY/mLeEJCRGXDS/nYS
DF/ULL0VSyUB4Co8Ztai/5pN1CA60qpA7TpXUl0Y0S+9kv35BFeVVAG2Pbkl7eMuENCFJPC6oWCQ
X4JL+wJ+sQ2RXvhXLBt+i8PruFPXBi7MWjuUYLmcDl0YcSpOEoZG+Vzuym8SVEjeY8TZt1nGlWEs
wVnnRTev+IGMraKa0uHOQrYfpCSyv4gSRGJMmtxCvsD2V2c42UzFgZYA8XR2F/9AxHkO18UZ9K9e
Y5srUnZhcwYT9oKdyrz+JTlUxrocObt4Dcbs6ZcIWCLCHqGghBOR4hsNQkXqIBqZ9fAP83+Krd1l
hoxquE9kH6zeZLECw5ZErI1ABqW9+26zHzLsR3GNcI3z4BiuoWSFjZzS+UDvF+P2cRlyNYQnAOfW
wWlR8+5HGunTQrLMkQgyh03ELDnqCFY3tFGUCjF/JHQi5I6Rx2BGlDSYT/w+swAzv9JoCXIrsq/b
wWbcDzQNmBhZVbrj5v3gp2ukt9ry3vZozY9f0XKhN6zKUgmlSS4Odol8g4uX+DdOCBVQtqQdJwXP
pEdQvPi4Mr1EhxYCSbZHGdhDXAWJy9p9O8K5vDN4TypPjhkTz6OoPWlNIMzzklJ440gVpDvK4K72
uVXLLAgGXjXPx2PVyPiIbZ9SRrAisJL+D78F8GskQJ/dbUHecLyYUiWJULcoalY58ARhiqXL5aSg
qV0E8tPQMGBxVsyYiMeNJ036vJYFS+PdmihBJcZNsEyjdjVMO7XkDC++XIs5IaoljmoBOifAMdxo
v5aUzwfcg9qi92ZhPhJmF/B3eXUk4MSJPYtgjps4/L3bloxTZC2/tmQ0ete83L2L5D2BKSIdteSm
vMXtJPAEkeBVUgucBxnOoDL1FPdj9a05SespwK1eUN64/IXTtHmcrlyNzZuF/rbDwxaO3Ujr2xlb
WnAGCiiMvksI6sSTjTN6UUlAuTiqi9GxkHQi7JSsyZ0NAU9ExRLnzYK9kcl34Dlc+zEa0yK/fkgL
XCWg4UpoTnu/iH37mCrk7qCfdy0BYHjzwbYstgk7sMwdD39RZliD4qRnSlQUcqfbv8FfxKR6coeG
zAhfOKB73R6G6vcmjIrdOcu1hRw8uO4uWvOtcFsVj9lxiqg63Cne/un2u9gmwzC0PFbQPmfIWfJ4
wgjiq7EcpFQk8ONyDQzO+L2PCADjEVjAFyJztzXHtjcU/t1golZK1cm5Obs8oXuBpfxKVU2SlJDG
+pWNhfw+g08SfZz5nZXE6npy/4RrnIMq5zyK6Pk2wUM4o0PAia8A+nV8YaX6fz2PUU4kC/I9GE83
ipa5hF8XQb6iOx7bWtaX0g47yqGg11Vz0MP6wLA4HDw+u9bTm6ol6fnEJo9/6icR4o64uWp75h6i
5svwVipWgOABqPnZQnxAcF+Y5URPgyoU4vTakuecbpwgVqbbTwfMBUvpl/j4gL2SB3M9xYeraYKM
14YzHrJ2gpb7orNykjrh74heiQuogq402UNZs1y39y0U98vkHePnKjAE6GouZ+xctgPkiW65br4+
MYTRwWCUBdRMS1X7qcHDRbMl/PJ+la4/sBIxfGkCx/9364Z2jauf97yly5hYuwSdABxvS8XPl4ig
tLmVRVo52hsuq/Hlqmol7oPQyvMwAwTWGClbwSqEjCrfjdrMgCOrw8QtRfjq7fUYwePMAgQooSp6
eo3VHEEv4HuuJ4iJDURgF2/SJj1Jn9+cjUiEPxoHioS5agxLlSxaKruXRD+3t3kiCOcvuzBNCuUe
+H0n3Jt/xpp1EU/M6shh/GqeYR/l2vJP1NuOq5+cllgqG+atl4b/OwUX1aN30XdcP8fqlQnicxJS
VZnjxYsrxCX8CnJbqeysrX7njtkxr8ZuJhlu19cNIGzrjPDBlukALsKQkfx8rX5jWvI367qACFbQ
oCtDk/mJwHHai1LsGrav2SifcYn3SlqK0wanYX5S5lqZjrdeLuEmzQSI1Z8U9RrhcsdR/o0mFPny
hVvUlmZhLUu/CDVzJL7npgawqt8fuxqp68rvVh0lLRoQ0zdD1EDSPLDzIo1JhFo0CSLHDL5JSZRx
McvkuiNALq9tByTPr0vIDn77ZYYubPe0O+iqH+B1N09qawVqww0iwOSxGJHJAJzYdUmVhbhTYq5X
9WwiLcFHoPFF1g/mBfxhiW7MabZ0AVa6eISbW+ib11VcWnqeV/OMQpcuUFcJSQGuADMYXcZzwZ9A
17Bj34qDNb7sD1tCGDPE0B5HYAZFXJrUpCDxGaavquEPzG62lVOvbP6FJuWNNU+rWyiFGdqpAFw/
DKrjW4uy7zU60pa3B15q+nHndkkPW600jsIYm2K7AH1M76jRgU+HMDxKHXo1vcaR1c6bkToJjzMV
dj40+x4e2bfLZiaEiSdToOGxIWfFJ7R9VOU6vm3kDr6CQYYyuLmLcuxlKqle74w4lZeFFxG6sHN+
MVuEUHoqzOcIcswwH4Ul1gy1M1D8ssSQ0FT1AvX/Qk++UpBmREnJ2jpBQO8ONg6qB95m6l4R7JCO
c38ziX8JiW9s4Ubq1BS9bu2xz9oQQBnj+LWITHCMTuJmpZWUk/WUnu4+6L/tQ4/umFp2cC5mzaso
uBoVkO0z5ENc1kDVd31I72Dr/Eh0UBn5B1yNd28m/c+0IgDMEz4fAFt7jVyWSi335PaWt2eY5gIj
HCU+wZ1uHz5K/yzJbhPkQvJBSrLwE/I13sdlMHMLeULIrPAOJ1e1M52xHkTWjljy2VyDvOLiV5Fs
ysXkDeo+Mqbq3n2Hs4R1Q9LDVVhrWhheoLHbzAabdojXOxbJrS6cN4N+dNYNlx8JOvAgpUzKkxKI
TqKAm0IdVb2DRcNrw05sHaNUn6odfEbCYn3cmunrYyT/7u7fpcQnrxt8GqDgGgkU612exTI1wZL4
hikcGM6zNQ2Am7Cb4lR8y8O668RW7ztd9Zis9Z+2vlSz3+RU5UtVYiRO+sOXA8+XbJRdXDviRh8V
HTcKFk5Pap3wIx3m3XraBIfZcShNFGKPZzveEN+amsTZ3Hxzk+PW3igAIN4/p+rZglo4J7RVS0VZ
a0UkiLXQPNAn173W9B4q/0nqFFaAXhypmOEWVuxTCIKhdLvv4Uk2OkorJINAb3GgkRYhzzvQtdoQ
mE4Akh5oTqU8lLaA3I2dUx9h5csL/WXZkjQjImSdy8rCMm1iH4ZZ3Az5NHRBQh/lCw4Yhyi+Ox/A
Va0bY2y0697cgtQduIj5dnfMBTmW3OmGISUh9G+k3wCUUnb6z674jkXOGFjntdq/bJ7MWvuYbiME
4bBI9ufPBIm1qGFv6FMjAmGfMnKil57uAGhHm11EJgqlUNYo2B4RkcmAkDxYKwAziAs61Ol6WpDY
wrmZrpfRd1uARS8fRmxu4zVt1WYY31eG01WIV+6k85MtXmZFJZ5+w3h9B5ZlFwcmGxOdcKiEh7LB
y1cFqYZXtt1xeGtpEsZDUsourZvE/yAf94lCQD5YA6/WB7x2bQBqzvHNrMr+M0XJPKEuBrTCMZHJ
4WwRtBJZWZ08NJAcHX2xF8qzBzgbP1Mo9JTd2kAYTqFlEdFS3KeI2M1FZz9DdpNG/R4xGhUzTu7j
icS7yN9UJgvgzwAtJA38QAT6kgaP1neHtq0DAxv1LvUewXw2bkvDq7Hb/M5ziwA3IdDkXw7hRCgu
g82mz5wmUQuKYKRHM/Y/PVZW+CA9yy51U0PVfHJk/yDV0djWt1BzCBpGZZp7getDkSGfyEH8qCtK
gHIiVUU2pzhMWfueHGo5066aSv2Ni0IX/HVxURdnLj4R59GjL5fzEmGR8jGD6GkpolOYCEABECG6
qdir4vKB18yq3CEQk8POqDoxFnAfuWLQkPwbpxZi8QkRZSQ5wXoiuiGB3/RL3GizDcj0zkOJR+Vf
zt9KcJDmWUxMF+Uc5KS8c3VLt4TAbCQpT7nbhoQf0w3X24UWeFjrGREb4h1nH+bwI8j44P/0C3W7
wr5LtJSsNl7VN2gj7QJCsjanQ0wzddIm3gqnDYEyM1fsf0duhZ9s+4Hwpgl6HRPVy1agabOR9cAP
LTMKZM8oHlAPpIlSaORUuBRc0I8LX4WZuLcSoUuuNqNneOOqC0v1E2umwGh16wnzRntJ+T7RGXcG
VbHirKqAdp3OPoisd9Ea2VYgR3rPboGRSfY4PW/hnFJdqSwq6/gLEPz9c3Thj+Bt9fCP5Hn4O/j7
840cJy3DcuPjxb55ZmukiZgVo5H+fB3WVkBra8IT804NJk8udVmJWU6VweVr7DybhjXHSjXfAbt9
DXYtt4QB/OOzPYHHKNODPKxcDi+V0mcvJcxnEvIiouOxR95+c7N1GcOGGY6mUzjV7r1JGL/wRwaw
Aiy+O0A4AznedxSVMFvCZaVq+VkVPbuK3muQSo7L6nDCsu8CbAZbRmccXbqUGgrgo8VhYjhKX/8y
h3GVBqkTphC0ljbfnJYhsgqTl9ebqbKcFFWQgA9Iqmu+2nrX4coSSX4aFeb5fpwXqI3lM9Hgd4P2
iRfeWXSihsaW3LMJCdvvr7mariqBXBA5ivFPvq3qpLEVb6QPJGLX27fk+6oZZhG8z+jAHYZQs1rD
lwYTQrDw3TcAoPbygJhEvKCsTea1MjT0x4KJGJ3iFyqJ0Q3i27gA9MuZJvCYD5V4Q7lSr2R25maz
TbDzuFLY9V1PJ9gqEukZA5+VG4lo0/Icnfmoub4pg2TaKa/uDkNjwnABMQCpwDZKK9j/g8shYaIF
1gcavv6BV0p+hiYbXxVrmddS53c6qB8EZrKN2QPtBKK810wvxtkUviDES3YTv3o9V/aythNrhx8X
9cnpuYMPOcs8qWE6HIL/R73wc1wKyDXW6DCwW/Gez/GDQmgwxDbine9P9WKbQpO7+rChL0a8sfkF
bv4Qrm7325kP6mTJiAS76M7flreo71sbDcU3u72A9r4rvRhrOVsgIxND2jwXlS1oKpYOirQ0E1tD
oOSzmdG9NKJ2iFuLQ0FufJSrWuR9VFHbd+Q4iyJHoJJrmgLayEmMrf918jrjVDv17PxX1rpKEsZn
GM9jF5qWAqHbsIRaleTMIJ/4q5IcZFPTzbMulMX+F4+yGTKqXJ2F7K2IwuzeUVMtK4Ac4uNntZ1R
xTUjhGwqhFZvchzSszukQQfRh4ooob4Alqii6BOvU98VCV9431Qb8BDtH4AbIP7y7v31tvx8Gr49
sBE8GF7Udfio03ul5UDy3jtYz4Hyaa5E5SbFSLYZmd9GTvBGg8LsjLPxydprEwZ6ms9AX+gmMhz/
mXKX+e+7SI3cPXPEs628xWJSfkGWjnq7ln1g671yIB115kOC8MYYlJ6pcymlrMlPq9LectQmaiXx
njrgOwE8Aa/PX5vOjqYh3vANN+C4BtmeOZ2FrJEk8vWeZ3FQnpquMqwt0PEvx7GiqEr8PSY4jv0E
yqhJDPm4SdHUMJ/98FwNDr/XmTlh4aQ7Sieu1XpKzMWqpbXjKRoE81oKlS9QtxdkdKX+oUVCEvlp
T72eb0FjVfBXmyHgltM1VJHkk4naL3gmO2EpQymfNdd5VUT2ZTQS+Pph9TJ9Thl1aUOtnRpMEPvZ
UekYWZCQmAc7RG3CIiyuJ4nFP0j9mVSOXmehQxEhP6Jf927UWlENyhO4jwTCgpOr+D7NwpFzGmzH
tQd7IGxQYyWFQuD38t4E2K61saDw4YJdQMrcKeuzkLoyZUyj22yu1SH+FjZluN1EmZSMJqbMY++o
0hSyWMJN9b2ATX51kXB0CNKtgYSuYYtEC/ptmjAJ308uLpbG0PD2UKkEH40F8OQWavSZ7vTTZq75
vkCazx+PzvQ8lHOtaeLWu/CNtnWjeXTOyX8LfH2mKAFDIxXrQFULTfuIuJYB+h75yz5fpcun5Xj6
V0Svi87vzrab+H/rya13hFzIx9XXegr9QdJh/aG/YhO7GEx5Q4amQRJc2VQefQcEtARxDW4RLWHy
eumyydwEvXbQXU26vcpIOPAz3SPA0KtvnJl8n7WiK9/934YWcQkmGgCqWSei6T3i4wqigARzWSVw
gd9lc6Mf464ix+RT3Nk8/3FBuJ8696tP6mO8fQljFgnlHGSWm4FTF6A6FXKjGuc9g7FWfpWxnkxp
0XEYrTgMUm5l2/VjEwR7ctHvDpsKrdtZYeJ52Qr4rew5y6i/inmbwJKcl+ExxARPI5oQQFodoxpQ
eB+AQrjkoS0AzLM+n1LfQN5IxxkbupWglighl9vyBVj+mjCXB64HOyL6wZaOHFF5VP4n1xkRCtme
3uFim2SSLWxH2vbFkssZjqpA/9gkJEmgZkPXanDsGUj/gR50Iv7mtsnJlqWnESI+Yrvknft80fIv
iYvvwDWr2JQJ61++/8iGIsNmelTlmPL+pgx+xqbynkDrg1YYRvCEQiq81QqJ766MVkC2oAFymA4x
eGp9Pww+BOOMC3iOj/bZMcZ+gpin0JkPZB94oT1mRxqEZIO3BiOfPVSjMf45VoBKbA0XgNEtEeB8
akOVdPXbJ4a6J3mDPX03kU+75k4yVbKB89zbfDHcAW4WrDCN+zpL+/3EEg/Xq0ft6GDMpBeq1kYv
kqB0xZ2XcEbFWbz5XY/3t3rMUvpn9mFll/D/xce2l3m6XN2HSeay3jtLeASiOUSuJrwaQoNZ7/5S
PyjI2yJIoV/CtPjitwVQ69/BU9S4KhqarwPJNFgcLvUcJloNwBHXT5eqSupvmzEeKJm+j+WVKOta
MJh4IxsVPb+PiOvwJEZ6QRALpfNvxAlSXwdvawWkpwZhEU6PF8SPZFG6jZVrkIv1XHcoyQM7nm0+
20ZyyXDDzDHbHOvFnn2hivyppS368qCuqERVNSdms1OoLegGqoCNYHY+412ShVl+On9HIrtwVlMU
fmA27M8DqnKy7+JuweL7GvggC7zEZ4uJtdagh86Pb62F/3UQ7pyKZ4MhXK15gejbr8T8uYDYp19k
Ee3RQsbyxYn/TOBmQjpFowKQWdHws3cn3Rg8KFinG20CAv5iQ0FMzmsTxioQcQhCyYMxc5/wfNrE
PD8E2cZiZP797oNmFJSvUKQp7kaIdXFl0Br3D7z4RBX4eRLmE6dYsLWcXn10sSmORb0awIHBtmfY
ioYQUEQy/g9NY7094Y8DoSNi+J9nAy3KWivDODuQYpPTmXlKfQWj3kw2XUYIPXehh0AytrJfbPKF
kLqc0dW9XpmMUNv0fjtbEqa95IbdE6WJce6VpUOM/qoF6yV1OnzCHkP5BYGRVFkyfQSWEV/zBa1e
QCxtVwM4hXlPeq+kMs0Us8U6PTTtVHcVJ5X1+qlR64JutASsQxKYj1AYYrMFFebYEbcTfL2cmYT3
gjms5Rx9h44cV0c6Ly1uNlC/h/yu67o6mWD/72TfwLiAB43c42twf4qPsOCqKrHGCYo58gGuaR53
LUL/2uYRiKphLe1aq0Ydz9cN+jjdArgN8kKoh4YAtLoVBjhNe0LuEYXRBbhjTTI1/+MyK98ch8Kj
uhLGTFzUpzNx2NG69tNeUc5C4CoIPzPLuUAyEOd+dxjcLQM18OsTLRr8FXuNMr1xRPoJFTnSSJ3i
dGEVV/cOJC0CUQqn/36iqkrN1LO/I+VpTKTcF5ZMyyFa3miTF2Qa/fGY9uzMkfqpsQrrRhuBq7Ag
z+szdz1cXOGXWvEDlFB76Ks7uKH6W5wZpHx1uHN9NhDpxQ+hrmdYyP27GcJ5RdPyLzQZDuqtHQia
wp1zUuljDj7UNh50DY9y7mfcwU6GwB7qI1edTW54tzEzKqE9hXXdNyoQv+hEmfek+02SXvapkpkh
G23sXAsUpS5/0vdPRPywa5xU+yGvqtnIILy4XBtCR2k9tcNTvpnTS4lAx9codpqrvCdEZUbNM+nY
QYJtCE+bNze3bnHWwW4tfgE8v85VSYwrRG0nl04k8hWeJidn8PrMb2UZtyGGxSGawvFx4YxEzSUy
GpCVWiphLEnlIIU61ioEASWfRt13cEFO7l2XFvwGUBxtF9sGZvlp8a6KLPUuUFjBy9zimpClLdEV
0bHCEhW1DOxX4GYUiUDqhHyPJjv6NVdgTlvL7yBcJnFVlp5IBANhYqN1zRBSFul+uNK5HwVDg1Y+
S/wbtc0CofLWWy9hW2AeVmxKcPHMOBJvQlIaNncbBHKGn0DIZhNGlbhULMG9ReZKeexKbb7mKDBk
/uxFudkPQMO6zXkjzjow/gUnsFhlFkKAXI54ObngHxs+CVOETyGhGLgnD3eF0rwKyFLpz2EqvtmQ
yTOmiJ1zIxRmkSKn/RmRVX4ChG5L38lV5/QnD2cIRif9H4JRBGLOxHqOEtopWfCRmWvaBqD+cCKV
uLtOsx+VGscr370hJ+LZY3G3aC/9krFRa37RIwSM4IfiiA2KhPR/ZqC+eS6seGaObZoCC2A89/Yg
2pqbblI1ByOYMMAzg2jVQdqCXV3VVDXOfc9+G+3F2tUxuNwxsoP1eDIzxocUzmdUmXwnD5oybB3F
fHzSGNKWnJpd37WYob6UK8MJOD+6CFfeIgKFmKAHFOK11NEzVgU1K2ExnnZ+MywEvFm6h3OB4vlR
8ols0b4BwR7pGIWuxnf6NBzwtRVBbookEX5xielGw4T2Wi3f/y6slXNZUQ9Bs6OtoBqyMqZZtyqN
w02ZToecNv/37Qx8DWrRoj1Ol5ZoWnEZ+cMPCVpkKY9/8/y6xwQD7UYrxh0mj1fsr8HWLiredzZg
ndEESGaUyFUuT56FXutn3mkZWgS6iXu2wxupktB/DBDAZvVCY3MJIYm+lzzrOtHg/WkRCPP73dVi
uiivN7q1qI+E9qLXBtSiDOJ2jaXZ3fKpPUnFrmHI6jHXP8k5I4y4ySh/XimOijjQVmMtOPeMKKQa
MRLZZwTTCU9OrYrjmb5t5fX6ap3b6XK7i5mOL+qEtrL0M2wyq12qzvqzrJDrRfWEwIJzj8Pkglgg
BMxWVcTbbeA0KtsAVdg/zubjN7Zp/U4IPTZrgjpV0TAjB1SpcE6Fil0SY/ev+iSyzMzJ/lJzDMu8
EUoyQrZmRvYvllFszUE76RztwWF44dyyCKZNLG2L5KtYON3u/D6p1D8eUxMDS5WtVtcTYnVLezNY
1PCqZEmgIncNhVtkel8FEm92Nqtc/AtRuSq51uWZSoleEDGYAjp4r1K0bGFdJAQSU8gl6La6Kqvl
2qutloARrenpl9UcWOlrnIafEt4hepEZllfnCUb4SQ57EyC2ag7Or+CpqRlLyvbBZRpga/CvsVPQ
ETyrfcw6vNGklZY6s1Mef8k4+W5sEVgjq+rsIQVL6JGdHjjS1IX8WXR8a83KHq1TpYrtAdqPmV5M
7SHad4XlK5A1lqQsPQ5KbnAlpQ+mwIHI5fF9bWsUd+sd6TGz3JIrCQxcHdTeJWrhy95Mvq5o0sbM
0ocjofAMvZZw/+I8RXhc2HgLPL46tELeSn/SL8NS8dFA0AmHCYCJhvZjRx5kxRPGZztughdDkvTI
jEGwMPlr6Gh9F6JRs42Hc5X23BhkaGhjFDQSFJaZv03L5tlYpM5guZxfqAST/KXhAVmOZpxUw72H
6ZIgK5CMJwiUO3WRqQWWpFrAKE9Wqhl69GWy/OXRnlq+tqrQMorvB3ztYRwsDeFK+W96zeHBbmIO
X5NBwzJjxIZ6Q+dE1fWdgaS4c76Oge6uWl8BW85L89oMu9zj1k6aJisEliP8GpXKTZVyAWEhvMi3
FipLfSsyUm6+XZN20omATGCVNgHb8rge4DrXSqQDMaRdW/CcbO3suyksrcXW4uus/yolWabDkXlY
Wy48N9fDrieQjosBGzLFlAROFr18xClDZ9jg6i8M48RDlfrE6c9L0h/qlmHyx/ig683UCiikaN6T
dxwE/ZcdLEKlfwVRc2zZbkkFfc97joQ/RKXqWuU1fHO6GfB1ekDYvNynTpGzReu+jSO88YUGFavu
9+z6sQK+SumiSpAPyA84PNn8Jwb44y64U+O5TZLHIAzgBS04xLwKFpNgeGemJi4E9kQ/izMzfn/h
PjldqPWdLTcWXa7Z7h2FLUEgX1b6T8bTLvfYANmjIsdzQny894i+N+3aaOOlLnb4a00WVpqa0D4U
kAzw8+8nmQgEf/PJEnS640ovtz58CX9+WsaZqAuLuyLSaS0DfDZqKA8FHCDmSXXNc+OW/LNwGdBy
n2Mjh5PDTL2huPpQLmxtS9pX2IjXYbSjJq5GJ4lokVszlyCQ804RyseCfiVAsivKOZYLCPPytZ6P
+1CCfBeq0jIukhRK7TRPgvYq47BD4WySInj+Re6KQu8kiTSX0TDB3x6H0Zj/46/9Ww/IvDe/EjUu
zthA6M7dBY3GM8lf2v3b/Kih/EJdyWFCDN6Y6y2WqTnpo1NeXvgSQsisuvu+peZjruXiKhNEVYx4
JdaO0doAIdJipPZA0W88B7UKInvViBeFABSqJnkeU2WdeXizzdIok0gUym2aMrRLtqlDOdWJlXqJ
cCVzJh1yEPsRrvQnXPDCMaYbLWC+4zYgYBuIW1eSM9JibO69GzGbLX2EdvcVfOZygCtHg0vhDBX8
0KPFNWMb27DGdgIPvoVG5MsANY4vJY8UJLs6/SgIlLmWP3quIx0ROB9rAVBp9+0sfZv7cXLZVzSW
DcPLuSPIDS4Eumj9WQENLVBAzIAU8qJLIDhjG+F7/91DDBJgUoORZLfSz4Wi9gWbxmfDUQYiyQ1P
RCLUhl0+zAbLEbSWd/TGH3CzS6s+s75Y4c+liV9UWLBBmgCyflhtaZwogKFeeabcZwsWp3hEZmS/
5txIE/Sutp2gVpdKeRF3UqoctVoHxI3bziEvkFQxcJzjLt67MAPn34/o5oUSeEaaWvq2zYLQC1ee
KnevUgPaQlDJocy+OPooc07EPTIjffgT4KluSUwkTXFq1sta23+XSvTwfUPXp8SieyNI8kb6SdPk
lvZbeY6eQRYufPE15V8WfzMu5LTQJsmoQsB6wZj7IOt6oVC3aVO0N9KtYtGiYheisdN/W5sCPHcq
Xb8AmYecWFkW4UAGMUC+XNQNGvbrgo3ckTdAOj+QpjZq5UYC1WIQBocMiHUU/tPLI1JZ3trbC0JO
7u7XliWAUEvPhGOHbLUBlmpd9pTCB0EhGrCiA5jQXWuwT9JNWLTw7qXUL1rXyIau4aTVAnzdUhbJ
dZlFMsisj0dbJU+EVTUQu4nnrYXoRuWlmrzYJrgBEnUU+eRmhosieqep5QOWlUKTooMjN0vF4GcM
noHxaoB6EgNYRUlA/VJbRfhdDveHwQfIZG28tP68OpqAkUjNA37/fFV3FhK1rXzJBkVl2ptf94Zi
wQiUiIjZ8Iz9gnBAgk7zdTO826u1FIKUXwbQ2UX7UvK/jh+FyyBj/ZD/ZBUesuxWxIR+Mw7/Ywkp
qgaa7qznLFDxJ6ehIiKlUqCs/y1zvVnfqYi7ipD0Gz7uxDspi+C49sAlpIoNMiUEaVLi5fON1ubN
T2TmtlHOJXfmUqAcYIeEpw7NDPNRNM6t2Qmph2kfiRBUmvUBRiz98L4HjYAzpI4ZSgPxvhASJ0BA
6PsWKKeDQW8e6MHlBsQ8EKbnPwxNWEK+8Zq0Vo7tDScWGpLXIEzbx5u1I/TDeZVID5OCAUUU8hqJ
St9jDkPBJ/zq6gUDA2G192xbaDvdaDtLOcRIgpAvelGt0pvOMRHT0Vy+8iMldbjcWkSy0WQpKoPj
ibZnojGiwYm6t+Q7XekVErhQqrTcroGiLjtDubArKg1cppdAysv43dzmu7KTAtD6yPnuJBxU/1yH
GlYSTPcckK/VEKL9qfyW2swmWauogm6+ZSGd/nVsQbT2TtEhJ3TBiHajU7nDP0lAPQcDKe3lQMu6
y6SjLTNuClvvtsj4q5xYgw+bQv8SgqqyBfZjwlha58r7SgfkX8TYJQIKZbPfmyd9B+lCGFgyLHwi
1E036wlSARxNGsU35dCEO/Za+UdBab3vBYiwdZQ5+xEQoulaQZF0mvjwSHZWuNRn7azWifkBUdEB
wvv1XXkEufB8akayTHv64KMjs8dtwWMLEPsGULhXTvoruBmP5RvRktfOL0TtXUiaM4Y8BT0wK1oi
dz+5KX1R6+PPWdGnTW0/2BMUwr4/QzrHoBWPq3XBiM+JgRzBiAnNimBkgxW6fs/sK8C7TKfC0xvD
suAuA2VzHcqxt3LX389gDygROQk3g1jnSTailL5rY7r0quzF6FnehJK/v6O+CfPsys7LV9gN6zpS
TJVfuYpehXRvTEieiCgHEFKvGB1mTErf542dVraFiapIXF562D6K3ywe57qGsEICpReSz2Y4iQBB
QHUs2FxEq68mhIupD7l2cCbwrkxthuH3DtcmEraYqXnblidZR+QODywCBnHJo+quo+qQd6QoaJu6
OC5zmIqHgQyiiKSOWjj3NZs4LAsAUWvA8JOubm9jrvdutDrqiojN6T4nQ16eKPO+aStO5M6nSgJv
pgdxy4MplZXl1SL+vWeKvTMNnd2zuM7D+dWUDDosNI66WU7lCoP5XqtbOTi9mi/fZduToJdRryfN
CGtUpCLZsQLNdkO1WtpqP2DAKfYnV+/S7N651o7aYMp6urdZGRwEm/gMIynhftLMKp7HKyrxGwhj
Nqyasg0lmHUtAFPeUz1p0PXezOJz2KyfcNz4O7HrHiV7ljOiq7MyLcLCyGt3VyDLKaU/enQSEX0Q
1eLQQ8zLy9CS3xzsaRxhZYFcnL3eaG+Qz8TA9lohaYea51Xs2/p0eLH0Dpi4Q/LSJsdN46BnLiZZ
/48KBq0x1uKA+5kKj7YDm8wpk/s7jJqV05uOD4UlWO6rLk1DWwQm3U/q3mxjHqpbB78xUd++Wl9q
vtJEzNm95mGCh/d+SvxNs+7moudeXI16cnroiM+t0S1BbRhVc+RXSAlZmCufhS90ci4jE9ZbHNFW
PLxYnuMj8NsMdJJ/5rbojoYmZ+rSnP42uO9rIuVWHSjtFHUgJGjqxXNZKXBkA8WCCz1ubm3OfC+D
AKHTIfg8m3vuV0zNF+3SP+na5nkGD+uBliM5YXS7HjMLLoOs65jDKePdYsdEpGGPUTEV/taAhqh0
F2Bin7j2NqB5DrZSOcBC3maIv5iTzxDwOLrV2T73YASchn2Ey4/afExWBeagTqHh7wGwL+d8lNOz
T2H0v+i3cyv7YXV7IzbGEn5JNkshpG7zrJKEbJqdkY+BI2BOM/FG/heD7PCC6D1ZJSX0pzuD6GsI
+mRsh4M7psLPNUC2Oqv21z3IL5rf0oUBIfPec57DY9p8rgCMyl6fbytemWCEyJcvaHuYtbEej/Ax
qgO3hBfcGeJ6pSSYWe7uiItRTC9RMJSTmn0xJwz6Sj37qPM8znRc3MxOZ+uRt4n3jwN+qUtTUSPw
us576BPSgGfo4ZjXB3FO04aa377TB3Debk85TuoPhAd9CYjGFp1dThLecp19i4jLNDEU/NSb7rql
8VtQP5VhjXRx6m/p51RU5LdX1YmMs0xZK8oQdPOta5u4EqPfYmRdQdarHnJSlo4HWF00IakRWi8Z
AqHUsOb/76A0ggpiHvKXCu/ThBsoFqTYiW/VUU8oB/WrPsDY+lWUM1UWu5QxQqemgOMiqSEskGgY
uZAQS+Lvrm4ht2P7SiYaSQAr5W4rgYQpYAjiwgbKBl4GTeMZgotSJTGtFVBk/wg3iHWDCyapieq3
JcaiHReX931umU3aCT0UTTI2A+eLcAwwvSpovCPU0mgL1JkdHcPukyOn/k+uFtI+QfPGCsVNA8Fh
SLX3w9AemwsKXB0Pkjv0jJTf79oBuMVLy0DSXWOqBowGfp+LWo0wTgJmAX66xkiGXdyRY9G/ZCAR
GDeph9d7FLKL9tyP8OGP/gi2IN75r/apvN2LLpzqp9qVc+tZ97hACfZFmlnp0x30IeiJMWkkQ0Ex
ZSDidhLBTC1yKX7LatJjliNZxeRi7bjT2Tg6SnGO1QwMfX+vxP2RM+cl4W6LIexSoCKMRhlvMxoT
X+eV53zINNloW+aohHq59Vy+7GmzkMevP52A5NipIjIo/V02dR4t+vuqXrPmfXwTiZgBvVNDmWjy
c8+EeFCT7KGDqeDuj41pvrgFfdwGmeqlJoZpdP0JwyX+ShmEJY/U5dJDETN4A0qiELXoo3VeadIM
d5ZJvJT6hg0iuiltLwlA3/ayM59T6G1w3Wmu8vEEcGrkQyxlYv9jw57wghusXRKlqJiv1uJpArE8
WsvUoGyw7D+/wvPzhszD4J+c9w+3HUtEq8PMyyG7dl/lx8J+Tk9kF7qlpzYjwwx18bxVVy3izQw+
fijo6tco/jXbybbTyRklt/aL3lMaN4rEB1ECqfJIfkCnpEBdEervXgifonvU8oSDtobW5iryTI7M
0aD/GxZrVYEBq3jV+C8G49Ol+v1UBqKXNonyppFx9X5KHIXoco74y7Ufy6jvcUWzCGLwjA4UPsTQ
XSrX1Kx7O8Kf/h3tfFGhgqpGV0qbHGYFT4EtO7CoN4mQ0INl9T1RGyoLlaWOnristTcMDF69OVQ8
Ge/vOqLjgVbaaiLFqLjwmS73pDxVh6mHaKMsJgWpsYbuM4ezdsXjwm2yyBCqjzBc/OYngt8nx/0O
nPo3ivS0lMsevDOxGMOmqSzK9V3cOMIuXozBvGk+wX+8CtfoLZYtnFfDccN6IqyC7kspB43cqZGy
pHJeo6JjFkrHZJgvN1PrEqUxL78YCzw3UJ9mhVgXEnLHX98l2k8VydkmYjcoPbuvr4PH+Hwy8WN/
KaviGhUSjd7FeD/BM9pPLK0lbR6skoB+aqzocMJ5yk2TMFFuRHu2kLU9dTGl+7fdAkFQhTGj+BzR
P+afwOWoAQDWnN2pX1GwyCxIkmtJKjuH+ay/H56iwNkWXdwQ2dwYtA1k7KBdJNsYw09Lzy6XCExc
uPASr5YGDY7W3o/6dBHT2CqeXhHqRWOQfjne+Ck8LCQxl+a3o84FBiErxisJsudXv2r44SMiDs5b
5GHyBH6slQBz/ZXTtnBTDLNtlOtxfdTieovPuKLukLIpR38JMQoU1OUPc1AQcmAAhVwmWq6klXPY
JHI3WYeht45S7Gwxna5UNNG64ezwh0oBPLqOE9cM6edQQs2mu22A9cVRRCU112acdGRmq1smJqGx
F99Co/n+2wtIzQYeuc+EKjUGmnVUfmwPgHTOjrz3asacQSvpqR+p84xN+qAkowl0oaUtivPzPfDk
HcXHdU/5fnWhPMpud/5b8Qb+CuIfXYtWjBeDZ/kmlkkOXCSl4fZG4LQCDP5fJnJXrl4ikLIOryVs
4yu5XE0lpfsTOyt/9RLIrStc8ET2IwDnsIMoR/lgJ9l0903Ch9l/GeW1JpJ3A/h29zDQZBrDAad/
alqOv7tLhO19T82sQPNEb9zBPEWfEzk2X1k7nQrRpg6UZu1BnXPLZXsMCdhfZ2f9zDz6tnbA33dp
lP1je6eX686iFm5CDwEB3anFx9gd16FklyES9Jd0im/F8TTnUPgRWXKlI5yO2kanNkEn7uKkB/gp
Glt4oqJesw9UowFFPDK1LzbxscB+fAj6u861+QUebPMmcYF8aeSBCO2Fv/o7kLHodJzjs+eY8yV4
C2OqekP3iZtIt+ZVTk+DOTCQjZsdc1RlwGzZyEWHFR1cqc+zn/74kfHWxXU3rEOljDWIYSc4HmVZ
Fvn1wF7J9PMj3VUIZlFDnkDstSjKkRL1/qahAN+Or74nGwbM9Mxpxqx78XUJsVrivny1pE1qyp3S
nhqWeTJjxcJdCghcN5uNW8lzJirReeZ+T9UrWR7iQ81Qt0taRLiCS2hNbrnQcBP1axQXNs6RPJiV
O5btxp1gQsAC/2n2Bo1QWxpjnlZZ0DPwbjdFlpoQXQTxDoB/1pSwOCRanbInkTdaK8fnHjt9tJFs
1ZM4EeNHIJWuJ60SPKjmfLamvbL81WnV19rxgw0AmLTPosg17L26yPaZR7tP3QMt4IAbG7VYkhDd
oKcDIjhuN9VrOa2urHEOI1WLa2GV24oATzb9IEP7PJKxncsV3erPDthbBK0EAcelkUL6l8g6TuKe
Qg5l3JZdllV9yNiVdmhu1cfeUivWO9Z+DHaihLfXzK6LkGyVLgJlSOg5eGMAjOAKja+DLyecX2vK
Pnyx6Tjo9AjhNHBKvhrhRoLVFCZ00X08l1f0MB69EdxUvosu1Xy6Xz08+GPaze0+5zf/hyYNyP/R
IaR4IlMBBSB+YHhpDaO+DSPeNlZ1PFBZNttrGLcpHNOD/+ckIzLKMi3Iae8eCEArliybUQm3EtC/
yZYa94KBOyy29ak5dpKZWCd9CPStthKT+eRCGmULY5fyxYUNUYmfYLKN8uuy/txNwpaQFoYpxT2X
mfNHK+fzOJUU5qG90XUXv+eIv+ZVwwIxud3WFo+g5WimbNbWMYMcMv3w2Or7IgeDiK455C76zaJK
xhP4+AuihE/8Tj0CuRG8b9y7pYbRx3VCiMJ21DrhNh6IITy4/k6jKQ0V5zqQFM1VGfYwh/Xi+XGm
O6QJMC2eIq4px180/kyc837t2QKe2y4QxAbPnrm73kxB3t5JvRkcp5CPNTg3WXE2vrHhUjAoQt+s
O5FKWxEzuUw0C4PTFoECg7GwTnjzyI3lXXUbnAD9xBJqe7LxCxXMmHrO8ZrTqSDBLi6ndiiXQJMl
wohNuupLXDfyaUfc96ynBFAqsiSPbEGn8YVdQm3N10c0kj9btMihAcj5WN7rV9h5SgucRYT3+73l
UL7AtbmPiNAwiMP0QDYUsSIMVDmNU1Ja1OC3VaKWD7Wg7Ea5J3eaWLJoWqnMCHrwdA7m5IgHNw+N
pFDjBAMUYrZInnqPEYVa14eDQI6hvMOPGDeXbsGWugbx+bssJoU0X5a1r08Aw1i7n8QW2T4dpegd
OCVQW+fH8jxqKguzLJcpLn4sf5hHy6nYGPPQXQAt+KQ4GwO309IccGN8JiVXZJTl/yGGNjeOV9ft
I2QILeNkPv7NNbDJZ1VUGDmQS3ONAkH+qlk57cByfqBLCMTZ8hH4wY79alDctcMa4iZGdQ8IEMom
IwwSKJgbXcrfZ4RkVp4XAALKEuEgWjGq6C9BNI0vfEgSKewg3kB+3Bi2+arLSmaYvO8vNawGmD2X
CpzHbOlco83AYGLX6oOAO3mR8MT3fOVvdpomSarSEhLkLZXvzOjyUX4y49FKRzKQIxiZJQOgbesd
xY49xF+lC9hOZgcuUDuunNodK3df09IeNe9NAc7TJiiR+Dj2Y+cy7bIZE2JlfprIsRkjwslqAzAK
GEprNuS9w5GRQ8xFW3l4CNTphNkXCMEqp2xfGNKhJ4rhXWxcYk+f28NrD1THmp+2T4nGOykNIKOf
Z4vChVyzlh77RYj2YdVLVSsuYs/PkpZzEDSDQK2P9w+J+5QTpudDlxfZZ3hbwzDF0KMYpDsEdkIS
wSc2yZSpoUtKeFgCTVIi978Vepws4xITrOLfzugOZCkHZuEBzrKF3DAxN9HuZLwtijEMS1hqg8jH
eZ1PxH9mwAvjYH6BMLldzNSM41IzXi9W/1gJBGyoxBFgYu+NzqqOjVDarlcYdknYykATylpFSVO6
m4xoy3xrAoXE442oKyuzrT7uIzQ5FB0ofRjMJYFiEboFfvf+c8+pIykl1j+PR/yS23Z2pmSiw+Fv
kfd9C5haY2cioRRAe+PqLYVKahZaw0YeXNZ0ddRJa/3d8pLj5VEHBYIoquljW8rhyOXdtxPvgY9M
5zhwSmRuc0RjZvT57Nx7QZxIKEQCtCZpuvr7s70L8Rvqzr0Y6QUvhRUi3MSLTJ7BC1giQGU+eKjX
HWssG8jpDwWfIRXOrLAutcGKmbr8t7BjHbw2zD9cWu5fzg7QRJc6plPG0XgQcFT7msjYaZHe5fzg
NTzZjtRrnb1TKvybpFqcekEQV0qvgkU61tStrjyhwTSBN3SccvfHlTEageSiaYJOU2M/mC4V1BM+
oxd8o6jujpfpGHw9I/cAn6JeOa1dNkC/CiguAWKDdeBLGE+V3C1gDOaE4QBF9FXsr9TDaqp8kSlP
pr/DaJQlw5zO37x+2qT+vL3C7FM4dKghQKFQzCsunMOwYu0bv0Z5rZlV3OGP+CEv6ll/EyZgIahS
Ttw75GhrScBNp1qqCjpvk54gp/CCJHDyEGDbMT3XGf1MW0ek6YpxAKPckqvxJ8r7wXC0R24R3NfH
Y0JNQWAKA/FemldSMD2TrMulQgKkv6H3Y4n6DM+3Agr/LBIFcLyEmwz+KTRjgfpB2QfrPAbbZ05j
K97eX3vj/kLFU4amBIoYmkbw8kmTyu2YLVBI400VZmxkNz/nkRShAS+pX9BC4TSEBC+kGtq0qqB0
JXNpKdB58pXJJfNBfKRQy6PS1N/OGbKCNUpID6v3TxvfVvwxlG7czSdw7qnlCzOSQ/4q1UH5wpDB
wdfJsCUAGDTOkEKqLHCpDVfbiangsBsc3VGXlIrBA7yQfe+l4G1fOVDApcBEQGhdwlkGfNKBdikg
LRQM8ykie2vz36DFMK0k/Wz90HLm+ZWHXrADOMZXD5IMYgkzNzsR9Gl3YTydnFB/0zoZbMH3/hUw
0Ac8d8j6e1oT2T7dmWcji04HuA690MBkwXbkISbYritD54GJ8i5mo1Mk1N9U2JTtWNriQ1SCNOy9
ke7UpE1ol+NPdQUZqGXi/jnUE1pkv4XllypQJuI3dTzGcPDRC5tWMY43dl2rPQ8WljEyiaD9nLNB
W6NJkBX9Pa1AwZjKKiUt/CIrng9szuRNF2N1TQ51WO7C/cyeEzqxlR32S7foBZqQXIEMDPFscaQw
Y64le/ThbiCilT0K6kdz3w9gSkb90NJZMGj1BuLEzn0K+sSRq5EoO8Bjz/LqNwwUvjUdZWjqfLoi
j+tvpUD5IeaiwOZkcgncFoop+ERMxcdGw81XoG7NT/+fzbncBIGh0pvuAQrm6oOSypjrcZVjWQ6H
1ZfYh1bSmYQ6BkNT38nUyU8ZdkgNa8GlHIzX86pRZPEXFGMlKgAk33HG0PPHBhZBia0SI2kwk7rx
YZcFLAso4zFikOE8pW/FFb37NgdfZo5HlFbF/yS6iBA6srzRyGlhC/cyyqI5B2YNmUG/T/lWaTrg
GiOmi6DJ+lZQUlp2DB6Dhy4tvBxz0EkcJkpHMxBunfyGGqH5zDC1N2jFNyiUXXzP2ioypTPsA4QF
DGTs86GdeOgZLGhYt1jRErVt0mhHGBGjixBBP0uae8g7YCFQnXxUUa84OOfAK7lc/hnhumWvOKju
RY9coZ3k+LzoaZsqnQ4erW1H/TnIzFq794hipuK4ZF5OqJeNozg46QgbXquCvjQ2ZOP28Q0VCSRj
eZAXHczhuifgYjQBoGLGJUsxABGKmjOnmeWdM5IVWQVMfH8mJ4kVMOv5CV/1e1JZv8nrarWagUp9
OKd9revPPhVixh+3PXqzjTRVvJvqS3cwRnyBavfGwa1tUMqE17eoogRfZA/pQQyaxKYifCDf0/bX
J3i2w66W7Xor4FwdRWWYa6yNDnluyJIdTUBKRB4Acy0C9KvX5PriO0fwH64zsE7QXeRAsYSjslH6
te6FQswVaiQblsVrPJvM+65oN7+/jruIM5iA5wxtTD3VrkCTZihAoniG0PspfWsJl73VPtGncUeg
jzDOuGI5b2X7K8o7EQci+xtE1NCuFXlVvYCJvd6vBkZS2tHR8j/nRZpTnF1gOVoemhed+tPdbiwT
4lc51kDePkPVKiK10rm9HLZJA03IRNCKiMftvcuTuWuoG+cLn73RDKzb66c9stz3cd7X934fLrAK
SwyiVNuvMH/EvUY/pNcdQsa1RlSSA8eznLnRGW78Gd6z3Ih5OL2CWrQdME7rtwFvrT7qkiupgPMJ
hUDlwQlxz4hHRxAJ4ASqrjhMMZT9/E39Ug2nE2AcMs+DALA7dReFEMjcv5Sb7PK3gPX0/Jw3CD8U
VgiZyuBlY0px1lzxZagit7C6IIHP5fdoWXKioaAL22F4+MuS5zyKT1++0vSII2NvutB4wdCmk0JV
OLV0hcw/68gx5sj4LD3Tcqpi+6A9qhK+cCv0f6l6waqEuK+j8pkKuvJBnK60KnTzVGtFq+3QCS4i
WbOp8gHz5Odq307Cwrjn1Q4eCfxMbJKQ59iNsxaaGM4PrZVh5ert1JNTUNLxSeaJrFpebA7pheM1
WL16BkW/363U7OqZhKKTFiM1jTW1bwhaQyX3lGe/A/4VBJFvT4a0/WWBD3w0bzpfhIdfzmTtgm+O
5Y3WQyQWcDazJfTOO09M4uqR2k9anTGNunxayKgp79xyL6iqa2VQEYB30lqY9t8W9JT6EV6CISQn
7whyBDoNHEgUT7ehGns89SwGnhXDbpcR7mYL4v60XqNwWAZUwjD/iy5SD3eo1HgRY2oxkDuU/NIk
ycQHWS4oQYFJElB1K1lVEIBkup6UDF5I7yITuivazU7iX4Cs0o0ED9/XI7Tvq9jyk1UTKBfM4hxz
bKyIVpyVvT+MdrtbQSi70eLuglGSZ4u+8an+eu6f+lO1fMZ0S2jGfBg52wsMID9KzRwfoTnhz30z
YQ2hrhHi8+6Tn1MO/pWJhYi2M1TjIkJCbwbIHdqOABv50t1wPLcpyq+KRuuSrQgJrtoUwxF4JT9z
90aUyfnS5G151mlv4DeGdMM7chsKwqdAK64RYULcmXVLzT9LF2kR8XOKZ/NhbxwyeM5zpehKuMfC
2yRIYmR2CqNBBbmwmbOj49Z8EqTr/oxNy3ak7PlIEGCV+BUNV41Cmv31Rl3UBjoKNos9C43wm+1g
xDtiDv1Dn1RKIXOtaVgr07yFs8JQI8GlDubF8gSLCzYGkXwh5Q8DnSEfaIsiJW4qj+HbX6k3hcqm
7y73PHIuOZ71BXl7eZoiL5Bsqrglo+bZkM3WepdVMf92recz0FALhLAMQX+HfZtTFy0JoivRiuDe
flPq36fUvufdbDS4L/nSZBGqlw7ys2H0528vJbUCCxI33vVy5qCXJFR47HNrOC/8jgCzW1CSRWVs
sXcZ1GPjFbSSPPyP48XCNLDq7oSdU84lsNEazgfUFETiOV6tIbriO6rtMeuIyhiHhH73tgyleXJt
/X2pIETTXc720tRkqaOrxAgGM4vg272ERFilsLMBgEfUhXIueSBnwx2jL6wfY3iXRSDB8366/AXo
alk+iaaC7FbfMxFjdmMzRiIUku+yRh4Bzl0oeUnWPRUa5hJoePqvI5PVnW10EO58bCnrsD/dnSOa
QQNBXPofCBNICtjRBsx7q3OXe9alwrOkxLbVCZaeqKzpntEra9Sjr2IZECD6NMisbkBIvNYULGta
RiOF4t4H6jeIBJKlNTtgQ+NlC3uk1VyFBaGkg+ug/z6ZhEN30sgVTV9Lv8drTVh8m23U/RUpoWu+
pg3QDNaiWIW9UUf/EW8ij9ulHInzEfbiNeHJWQLSTBRrYkJK5GQx9dKgWsYbE/xcw8UqP72imw/w
tTnqLVn+ICMnr0nzTMabx4AMugasADFBR0QBOd8wq6iBv1NNJkmvwZEuaJpIht5VMDAwI5Nd1RwZ
ap7pn+HlNfEDo2EZPyKZJpc0JWs1yFFmCdkQZlpZNlZcdK1I8BVzCvSPlAjovhNC/BH4PL+ub0aw
vFIHZjlS9Tx+vh6/WuBxUeRGPNZtxT8gZZYrYIMJGeRIhaKAYz573MmRLRwKYy52pJalEfhU0Buq
Kgmp5WCgOiUzsWYVi1PBNWL6pLfGa+igRStxJglGhIDOjUrYagUbxZIxVfEk8n1V1hjkiBgxHeF/
hGwGGpp9ml85yaGYLfbJOu0Ws+ykRRfq+b5WU8SYbH993ur94c7Ox4zxvA0mJb9Q5QaBsSGDkJKY
qZbgd5WB5MsqAnme+Qt7dRE61YgCpe/paZ0jTNiTxWv2m6u3roaO9X5KTyHyIL+RVuroVa6XeX/3
oSBck/ZmqaVzxUZOJGyl7CNRO0nnqA8NhZ6kG93KflUElERq8WPIijuRaLNOJkOR2CcQuwcShr0X
9KocokBMuGcNrYvMDRtC+nWmORco36O0rBjW1qgMonfrHrvdhHccapO8OYB/LiJt5Lqfc7gRlH/o
JS7WT9eLaKbiSHPymrAkdkxRMwgxLvoXFMFeesxF09GrlfgiNL38JtS0r8AapNWcMQRvbuW2dBPA
vHtC2GkynUhyv5+uvZXv+Y6dKxn2s/BG/AHhx3/t6CeniNvxVokCshCFShp0lx5MOXkIR3WhKK31
GSbvnOjCd6RAnc6WTtxvLguuKt7TW/wtDwPrc4nRu9n75ApyK53VleYt+UfSMfko3zWJDQvGgHcL
lX7dlVhz3i0KkpnU9PQT+KydU5s0cKI0EFqaDZFoHoOFVS1BXKO6xqKcfNP9zOLFV5ajioZ+Om5U
412V2/iOtgqYwCYu5rz0qh0wTaYtFd4ThufgscstxZ3jMUgprjfWUL6iq2P74WK71VN/FspvY1ku
EEtZwUMOV+jci1kAVfIyyJ8g5VhqoLCmLgt5JT4yQYqEFFLwqsNBRuJsranHzN4ETaY9MzArolF5
KH1/OlKtEJmYRnGmSv52BAfgtnvR7gYfhQsxGyxjPW8lU7UTR8gBwBFg30lTEg11BrClu9CGvSn5
EN+aaAF4MIoOLKtnYhW4TdiPJPbUPUHooU2r/raJ2dhiGbpowr/xum+MED+hPoNDqr7HRfCFHqPZ
4VYDCfEbPhZ6FvI2iRE7of869z47EMLK4v//2tfyn6sg6P/iqIt9RCHSZ8YU4hcoMTLu+PZxSCJA
etyuJEdoTVCpuI3UhNIwMw09RHU+tMA2056x/KbyDQVDNh0/ahdgrs+4DZpYUfHfJQ0c1qoqaUCq
6GdIfI7JIZ0jbWHrFxC5dqCUWSLRl0XwMV6S9P5PIPu6CAccIZ997o3lYN1jKOdmsX3dlEHa30Zf
m/pE/xBFo4OhjdtZtjmXwOJ5m+UZ++F8e/TjRDXAXvz4wqRMeyrGD4R2rXsfexEysHWEoEK5aypF
FTldyq1JIxUNWRDzrIt04WeSANqrnya33zwRT35HiCZuwWH5/JrGHnaLz+jwxVs7CEcHjQFqZLEk
sQcqfWxQTIX99/vMs3FRAYF/uzYJSrJl+VvRyGcU2rkOZzQptqWr2deryolv9vvyGXuGiQRM5Mj1
21LiHWuq26LiEmX7PMlJgy5wW68bzAKHTIC61AeC6YeaSinbtNaRYX5hDrAdVJPk+wYu/OBBe54o
6tREZBTWWz+FpTuS7HZ/MaCEyybmDx2u1U4xTCGtoupqRlXZt/5dQEAPHAzzM7RfkoGZX/HXwP6M
lHUq9h66vCyIAaqrH22nNhS49MJm4LNuPELourbU0Eut9OTotsKPliR4ae7asQlLOzFbpWYnS/rP
OqIzfkdzDuxK6/y31+V9hjvPCE01Iy7/5xIf1wHuBvkvykURpZbg80z7OQnJQ+kt1WKl/nPlg0jm
rHensYxIBvsXNrbf6qBym4dTMFF3j2DRNoTpba76KnGd5jdXVAo1raK9XiD20UMWBT16rwlI1ijz
wXqkZ0QlQNs5isrPxpzayyeZQDj0EYY0pE4C8fnwjIaneyGy714WQrC8ZGSXhSWBQ+TBJMU66CaT
gT8YzzSQJfBGvaUXtUE5K6E+pAVLOAuHPs9MToPVBqYfFiWQfTY7aparz9ifZO4RfZ4bBNtpPWlE
FDYKSqnLWPOp9qw96/2iFte0Nx76Ryv/TzT+ISbJNOF4T1HwYftw919NWLOOP4fukWal+LpW5IJM
ns0AT4vgctbCZI5W814dq58PIDcnPJCpBB7MeGOrvtuIlXLKd8YRvDt0ADnp8qARYogwFQbt2upe
oT7hMR5iAsSZ4mgFinjSXEfN/nwXKSI3btsS2n3lUX12aD0gzysEDsN0inamB7J0wXLvt7oixP+Q
FJf4Px8+Xzu8puQrFLBxJPDqGl6s2coAVzA7Jm4DiQP16jVHeAlkS/UD6Xko4BG29snU/FKEjK4U
o7pSLDSChRe1OOHYb3x97pksxppqeJi0zk3nh42BVelADpayS9NNfCY1xUt7oSWYe1k9Lmr9MIp7
EhPfJVKEeipyhgVdaTfBdKyRAEHwX69zjTN1Q+ufhjcvKtdf1hyoXoKyKPlljRrGE30kjLZYZS6E
e4mcgoOD5zw73bowwXan1WItQWQRfQ1BQZ8xsXSskanxOnE8xqX65feX6mR4kLvmYJdSBuPpExxI
CJD1XnrIEnFlTGn5vD+bSWZ/+XnQKrAc7cCqLalMjkPhfa7LANIDRODaX4l4TB6xlAN9HWaSmCdL
zVPl9678Njt/UMX8Uc7FDF/d5JHWrzejV3cF71OvgLDQsO45hQ6KJB6Kds/d/QODci0M3E591Y2k
hIO+NXU82xDJLPW3CnWb5UgEAxq5CWWETmjjfWMHtsmfhAF8l28N8tBjNHgWSSJbbPPW5LBpmCaw
ECvVsZMT3QfJWA2U97PxRYUb82M6S9wc/h6IJNYguTsFHrHOaz4WmBR9OytPq2GN5lAqyOJR7GDO
cBzQriBEB1Pc1lRaR1273UXA2fhpirQmVM973guMjKeHGCC/M58J3UWIeezYYaYHphX7IKauAlL6
i02J4agU3PmSHb7e2wZ+EOZosgZJ24OJv5ejfkM8e1km2Y99Zm2dHnnGgaqnCCxRdrSxeukOQB+X
77p5LRbvW0UVbf+Zb3r8GU03ic90cZHSnLukYOXSupzIKRZYqkkoqU4TBSp0FmBKvPwV2FRW3ytt
8uQuSJBtVa2ts1tb0Mm7rbfuefqeFMUIhrpf+UgqkZdpGweqXbM3DdzyW6F/pZxT00c1E8eMrLPF
wOQ45uXue0W9um6S257x69bbqlkJ+iOGNa4gv8FGccY4BVLDWoqI/tWlTasYjxO2S2B/aVkhsFqX
gPxtkjLYmfltu5GuOL8DKyU5/6bbBPCH9tXvZ9sVxFrBOrNlT/Zabq+pmyEZQ5W97ZvE1gCnoDFh
SiBfasmHsWLvMx/T5U4eGnfBd9LAqSZoGHUs6LIsIDL9x9l45e/HnKM2jqUbx3giOCYH1AxFrdSQ
7kDhV+YrbVgtEf2qnUe2IJCA+c5czWShwRMj01AaEcf4XIZnhG43txW0MohOAcj4peh0C6iO01we
Y7qLmyBWzd1KJAe6vIWvfK1VDEkx1P56ldNTTKyxG8GCwkuUKan2Lh2DQmutMome1XVB1wsab01S
rQv0kYF5flhrfXwkTIgLyHmNxNg8CljF3J61teWxuC2e/o72A9LILPMy75gE4lWgJ6TEeUNxMwUO
lbwsdAl/uSL5G1/dqSpxq/auKqpd1ovjWzspu3dvOoQtf17ASEBTWcQndZRL8u9A5mpKjHPI/+5M
NbN0ZG/ezBSOOzf6NWKdsak4tqOJh+n7HEYvSJnagskCXVElwnZyTXl7n5PxrzTcQd1vilqNmTod
bZzFTiTcIBA3AVXWrQU3PYA1IOGgcS3YWVfUCgUscB5V4shcWMsPqTDLbBe7PQIiTYuk1qEYMk3x
n5ttXCB08l8Z8RfMTnTE6Yw9zuSzQFoE7tCdHVgfTzDbp7WI6Ud7vMA4vfd25+36h/G7k6sd733J
AXVNx5r65cCyVnhtDNTTKw1fQBiIHkxDLAf3rRXNrXKL0BzLpTpqYwS88EDsVnMjEeU2nS5Qj5H0
63Z5Bhv7ixl2uGOCc8oClr+pEdxuZx7ycC2PMKwMyuwNoZd2vmQD3+sat6LOHuIxzYd9Belu8XqF
f6JH8kJeEnlhwy1Em/bvQIYMeSux1pssSxqpP74VsrH4zpmhmytFXFyaGeBVYGxvGwT4z9W8zOxC
fCuhaMGPbwQJ5hfb460gcE2O3PCa1Ny9Qp9kLTDJ5xPo64QOYVbIiv4mTFMo6hQvvmgNQkqXXn63
q1I7rzfaKQZSfX9k32RfWrdyFb/S/WIxjfkOuF3AYOKiijvd8AspbVnrJxfDzg7ESaNHj38adVa3
g9lJhgZpcqu3/qsgx9d6bZaMOcRBfoB3Uhq7QT4F4CIcDV+XprhXkHJECRk+zXhT7W/wgWzZLCXu
DttiTPR58X4awwBRU8zHOOnW0XQ+ggLxKwYS8qDCr1h/pVzPtLa7CE2c/SCJ4nkqO8EwbesiCa95
ksFl+RAQSBEaW6iqu3lO91c5sNFyjzjZT4LIVgRSbm6y23vFnl7RjMLdjwO2u14mn2PJq+DLuAHi
9G6BnW3/pBESK3JIFbVdridkhCSpkoaM+H5aaOCEEQIVUxw7dmY+ZYbLScFl5XyfIjDWs80+Q0Nq
/VHqyzkxzTBZlO27Icl/1mxsI0uKYPWk9KAhZkXIRKiaPt3DaqaJwHEs8+/L/RUO0cr73VMnF62G
+J4JSsvCR0pmhrzfw/XIyz83zQfymd2TOdoXh+s6WpB2VgAsksArlVvzaP3ZaNwVcRCvg/D/6vbr
xVm3zMf0Bl4ymR5KZziFSherDdVRbG5Mo4qkcukreyzxpV+4G3bZVjh2UPu71k0dhA5CO0ZbVOBg
Lc83y138oiOdOOZaUUyB2d+wZzzkKnpt1jh75PoYvfoWOzF9qZPOC9VbcWNPTHlFelA8Bu7Ul4Ys
NhGm+/csANLGOqJhbFeuOyiclGONPbVuvIG7GQZTar6PsifYnqqOiNXCk+JY4UNbec/VfJ5H8p2h
wui6JXbujMF+0ZPgnytkC6AOBa13faEJsTgB8g8ae2I6Xz9R3RU8/auYYa73S1ZeRi6pZv4sz7KR
Q3+UdVcB5mJAN/xATlssMgI9/dUVdJgOpHO/honyUxt7CGizoYlMqursBHlKkdIvhviFsphO8ZkB
ldgtfq1e0876rJ9xwo6G8ItIAgHDOM/m1Z8X2AkKUUHqne/GQunQXl1xu2t+bX/kpj22fwdDoLiQ
LHLvTUAphwqPOlZz6XKrdiqseqgyZNCwcx1BIt8mCVmyTD3EfUfPDQ2bcZEB4FfaUtcAsPtMy11d
Khlf7xjWpx7fsB/kzLNZphrv4icIs4EC+wt1zuCqacL2wx8aT0mRUiTc3I95hLlSLKjTaTHegWuj
9cfG4muWgPSmNq++p9vvc2Ee0a9PzLvtvzaO9RX7IvHBzC46Ut3B5ISe6FyQBENhihAyDJsCLOhG
odAVN+wL9Ck5QeAdNvF0cTJOL/QfRbznWjdpVSnypkNaKGHsRRFltOSx3OtNY0DU2HF9WD0tL+pd
4AdyRsZK4BRHSLGk1rD5oOcqsGreDdXP95o/b4TeDj9aKEQYNvqt+Rp5T/eHDrqSQ/zHbH5lj3AI
84ibDCoaOdrWpsFa8lFaeevnKT2p4Gega2eE6OUvOzZ5A0pYwEHnVbFS4pRTjMW1gRrqi/+6j8TP
pllMSIWyHBgqFXwdrxYPmEiNaXDa1T1kBJ1v9nuXsXGWMyvEqVkiNi2RakqDQo9jt0JEqK9xvoBq
H1M0iyWBb9mjr+CTSZVvDqiNjv/KetmVJpvPtB3Ptjlc2vtCG70i9hhh8p+xbgIG0DZTfUaWT/wP
HGOxfKmY544V8Ti/rEGrUD3ORbVr3jcE9N4GyeIjhYBj2avG9myhVhqn5Q+yQKT/Pcdh5IJCTbfH
ebyj1tjZyp/qocja+Bl4Hs8k0ttdwEgS3Zd38TkR5KT1IJ3RVj6yzpFG2gtwg7J0136rJdygzaiv
L6nxipm7F3VkZoILShb/yZfF+n3huJjLlDF4XA0r7SKsdjn+wSOpuV2xWftezQNUvk/NsD8Vgzpc
+yZiWB9pgDKiezf7dtGztQzQKp9k46QlmJhG63jXeRe2G8CegO5/QYtynBMa1oEgKII2L4RJuhro
dtQagGaZGMKm82aJG2xwiZYdWPjD9roA89W6XzB3E28LRJpMBv+sCS4LG4WQDbINRyCv35WpWbDK
APHJ7FY5MJ0nMXctTsUBbzFgSMgfu0jg1ZQ7HHenpUP0seCnThwAk+kG2Ul321hzwpXGTUE+dcQP
iyl49DVELy6AOnECUB4F0M33jMd2oYqSo8jHz2ZtMiSt/wDzGuicZrCWGLTQnL0zoVl5A81k+Vx8
brcJ0Oj9mlx4e4WhD5gESpfeM2YfW0oBJ3Ai+GYtkG/nxSDYCBecN23DbP/bSx/7piTuLWV4U49b
wW4iCVkUX+7ykkuqGcDAEhJ5p7l08g1WmqEd8QlpeSGQ120/8I2pgUJ5jllJNbwnx1tBwzPE4yAy
b5lTW58lNkggJ6P60e4lLULlW93Zf8+dkH5zwbPrI8x0IIcbcc0zGfERjpDKslFL2XOmZK45cj6M
HGCfkPU8OLIouDfrrK0GDc1bBozYl1W4UH8h18SKq1o5dGSAyj+ZB+Tm22XXOVV7Wr0vO88IMRRV
oEogsT0ZFqaFxkNGTFKUuGLl/X142oOWi7ydltyISR+NdKN6HHQNyYwq0CB/dsYi9mpWCQ+aOqs+
W8UtFQIffZh7njzI+9xPu8S2R4xYpS5P3+qDRc/R81qHTPB71tikDK/rb13ii7tq5DSdsGHjaORU
QqgdmqvwSz+5wz0qyaIw0rirFV4vgWNJUCcoZaVUVE2GgHddwq+GdQDpvcQ1tDrZfhjojsZNv+qS
SvVZvlv8QNevygfoqZm0SCkkMtZ1e0MVeWVag8194IupWNaP83e5WV2c+IV1qabAWc7kTsBQLvyf
k8FvQhSMIqc6KaK1xAPXMAicI1ooLG/SfqOPhdFA5rz3d/RpXcnlzpOKSUvN651aERm/HWLBdy1h
tZ59Hgv9LPwK2BkKpjaOjcQR/zvAcuov87wG/ZpTvy97nadEMBM/3H4tswNS1jsJEHJ6NRsb+TXU
qgoZqNXXmr5EzQDgF5HV7tBnLnALMt5gRidOd7PAGAusOoW9L6rjUP86WxAe2QiHXo5+4Dm8ajXR
SkiCTAN1XbL++mzd2nVVrWQ7a9GIPRgyyLQYtFFeUJI1ttGyfCRz+/CgrVyTQnJuzKVvb9bHPwi2
75sUtNOm/j6FBZHiilTrpaXTGgfWmv2Tr825LZSOGpzpdebH9fV/8t0wYumpk7oubBXigg9VGSSS
RjHFMYnZrJ7o52KSw6WDfydzbNUpo2RhiE2xYDgv41GtFQszx/zkdDZ/crm2y7Rqykaw2s0finm6
K3M15ZsDkpRgbivQO6W9CmV5FXXfpRKHbZ2ONoayOXcUbguloL5/OzefhGk6WheWwXhMYScLUFtj
WubioinF9LCz+8Nxx56we6NOxQtq8pJncnKw1oz9FyKBT5GB4QBDWNkaqQbR8oEFQ9AUCG4dF7Eb
7Vsc04DiQHD2/R/JJgWUxkQe2b53h6e0Xm/90xMq7rHszRPrN1XilW3X9MOR+Y5bx8kU8oMzXt71
piZed9nyoZZjN+Ld2T1WV8pct5oRkzrv8ZXAM3cxGzFoRprKdmpgmyvC6B2QzifvGsRgYpv29FsE
8PxLRLIvlOihx8PmudFVgCQlE7ooZtR9Sm7iujVpN7ND+pc0Horl+/kfPPCFcGCYu1YSIk0TzZO3
DDPhEbE9uikM5bOQxA/LzbHyquJbti0ATehWwawHHpGWGgKqWDAHrgMTxUegbB4cVlwAYH26+zCF
iKXGQc2F1UrfDTclTCth58wbaliOXWMttaHMXsL7wktXZDk2gIRDSbfUazQuQ8WbdE1BbIghAj7q
JURbOGCrkS7ThOaspQ64xbB/ewGQjN3X451FuUaPgLeiE5CWvQCY4lHekPZf/FHkHsCG820wWG7g
M7/rObrRj6gwD2hCCPaFhBeLAPpaTbMOn7g8F2ejtY33/HirTixK8CvJZnRAdcFIK8PxvD2BtD3m
ck+UsRf9Il1gnmlcPPeLuvcOnZqcOmMpth1JkwWS0+KofdlPj7+jwwmFqyC5y8VAFX5+uaKp1saX
wr9jj7LAR5LuB4c+eGVF0tvUC/GJd2xFRdhTVphrT4uuAHuOuGwoWFUKtI5jjdipICTD5OED9BcU
5aK5PpHOkFOaEe+adkF4sv94aWyLAEVp8DlnL2+Hx754Kzj+FIBB7eK5x8qpa2eJN+1QW1baWX3u
DGhqkQ5XBAe7BC76YT2uCeelGsxzpk9AmkGzMwxfxhp9+u9cr+bfBzL+sWt9wRAyL4O3PzrVa8V+
nVdly4ueFvbdXMD+EwlAdj5DseitEOgeTQnnIcXMn3kOa+jq8b2LUfGPJdbBGcRpOu9GuGuwcxRM
piCQny1B6b7eDtq2KXcKJTIXcQBEgVatMDVJMcKsYgA5vhJRq4Mh5j2nikRe+j9UZRDVy/HQMBuQ
9t5FmVkGs8W3tOy9sSn8Yb310+bCJNYD4ykqo+UEWfiYrK1/oPilJBIrVypr0O6ykzZ/qFh3pGnf
iEsBLB3/VdNSiv3fxCVYp/yIUsz/dkcY7kwYfb12KJSq7MYeDMM8b6KqykOAye3X0nE6KIGsr6xb
xDeczjP5HYRhIVvWsizTAxJrRqjIei+81T7c6YMlpEEiP6xMv8SX/3Y2W9PlnM27CTiS4jVYAly9
dz2nm4dHhrxNAfxlUhXa8uxG3D2bsaXPpH3GGso6ZtN4/jG3/UvcDZwx8RIwyCaib2UcsJhbBGtp
1PbxNNTXwjThqfcogIqA829OxVoHBs/l1TI22zDFFbNm6KvAkqQirWS9w+RNf1cm206I2FvyWT+z
3dNv6aVHEn1dbuTgFgFpKynRrH81JhRjtVMzKixYTuMCno5zW64rDVc4aM0N2szRk+Ij3XY47ee3
MjbOcpkQX40/E3x4hUYJEUb7WfkBduDQ7YaTa1PjweZM6zu6JmfB4GGb16EyxVkW7Mu7vB1+zWZ1
ki3a+B80X/iIxbTCpeU06G7vJ0LFNMT7z3r6BtPN/slNrKZpKrOZvolLOUzOLl1foXEWy6BwrjW1
/nuMGWMldeE7Jjp8SL/WVSJT+Z+d0Gl8vRA1c6iyiLlxlBbefSSR4P/QrAo6uMMfnD3+jVevakB5
WTyxxZjTAGtU/AVfevMXizOJxhTGpqPoQ6zX1YBaltH1axocg8hwFzwgrfoH9kTwxQFl5U1gvclS
9YgVN1R7b6jzpy4qXr8y2AtMXwjc/5h238zRZdPPSUU1ApG6JlMfWBu1vmtH9py/CxEf3HcZidR8
9+mRyG3unfnCEkc157es6abQy3r66dpI+RJc2xkjXClwmDRKj8OnSiTX6WryOXwakStR+TVCEU8Q
HDqP4gdgtcD8y/o3LvDZI0Xoa/34C5ormJxpAVkih7Qu/uADGCTSynrrEHaRJYSgy5WZPALGJ/PT
eaf7ukcTL3Em5OXyrEhxhlQqzKxwM+G9D71b9gJDxZAf1GutcIXksj8BFZ5ve6WvK6e3sympXP49
Wg0EJG92intMjreopd7rK3ic1u8Fj4joTLXkKqQ3KC3RHrj4t3FyfRotE7YK7rMOamxuMqnZuBzg
X26wZf6qkznRQu1OVh5n+FlvK9fQLVK4lB/Kt+xKtUoaUtpv7uhI/yQ6/rDTyhjrZSFowigwPXWz
DryuaHTRbNWquDSwT1/7++oxwDzEbbMZx8m8K3k3wafWZNfcMp55+JWAQ1PPBLLGVj41CqMSbe95
2TfsDvD6LC8s9035navAYQWwhcn8t4mJljBvQ11h03MVS9x+wIQvF82QaD0G0wS3phPKtLQX/Y4d
jXz4de6K7rMnothNa1s2bAoJWdli9GpQ4QKjDy9Iwc56KfLtavVon0PmkNtqVvKDl0eOiku0EoF7
/0v1vDDKpPHHDYfcNMnUyTl3Ts2MKu0B5U+numB1W/5s6TDZZuMZe84nLMQ+tbzqQzImbXr5Ya9w
tqDUNei5uZ6UwR/O28ZH8vsSABJ+mKEMmupbrchXFI1cOFHzFLBSCtHa3230IeZY4xZ/PwV+rkj8
38SnMGVn9300nJn2FJWU90vfqy5XXy6JDpJEMgXGQTpGFagY9eSjvl8PVo1oF9zdaqC5Xpk37FCV
2r6odjx3+/x2hcbmEepvakBm8bWZBFMAwtLLAKbDsszUZ1JNJzSuST2tuZ0cgX5Vopz28ne+ECRA
qRW3OkbxOxf2J0mswTHnpe76l2GJyt0ZYeW3cdc7Fr2pQd1yfzCEdsjztPF41UjZuhfcoWidg8Cr
HwEpV3RVOa3avPOBmdfdRZrJEWAksysxEsS/IJBm1nK7zgccGlaZS5eS67zTTsi6Na38AcZPzfBu
49DprH62uINvypZZPscczBfcBQHoD57vNJ4DfMi9jAjxfBu8WA+OTAU3EY/J8Fe/QrbJKQWXCEJK
MrvfGAYG/CoXEC57xA1j50qo+ojFlzQ2CJ/6db4wTNzU3qHuhjFe6aC9ypp3vB7TZ4kn09Ge0KG0
CDGor/3WopswCGWNFdyoYH3hJERYi6ItAClp8PZb/j//XxtX/kzdq8QaeZCvUoWIY0LZgsqWs+Ay
aVfh0hO34S8140caoxYEogc5skLA3Uit0NFIVQTi31VAwMmOoxx+9P0GOgyvxQWYrWn/M34M2kx6
d7h9jrXa6IZi/JiboVi9jSOrZRO7mKpIuFzEfQcP08xthKmcYkGSI6MkRP8X2dPJKSQ2xNFJpfVZ
kbh0AJzddpSz56tNkynMAenzJmR9X8jVJXY2lVb+Ex/9gjuNBzgz4Ch2G7WqSgW2inqfvFQTorsS
Joa3gb5urNwBxGiFLp7MjWbUyM2bGusBAmuV7K/lP0uVC3GBOK33BRK/Uz/pJGT6NIgYEnDS6sh4
gV/QDBC4iQX18MTdcNJvU91hRJ4/h5jxJdlkf6DFhxN6xqRjXcSrIMR/bkg6JBB2WjPn7g+0dmNr
SwZ8sdI3hpQc2XZHfl7mT1eNoh+0Ik0YZHbVStm06Cg94j6fmCwuyhGhKFqT1YV9jKPcFHI7RIMr
1XWKNn18PIcOTFexDjAwS+FOkCFhnHLqLNny67MIxtez71l/Fb1/MMqkOZD86DIvI4cZhersSNol
+UhJpGvTpZoBxd0FNupxsWCdlsfCrMWQFRafFl1w2bk6FFwGT+qxchiliI8bCv01bos1IQo43yWg
PKX5auRP2VkETYDR3j/O7XzaeHzWCRRgHIR1wGEDULYN6rNpy6vhN5ghquJwrma67uYsIq3DimBA
X1TeZKxHl3DB8Jp9Sw9QdKfkx7d4Alf6z+qoIKZUUiaKbyU3LWcInE2FMNKtHZAQkySIPGacpTWL
HDTMLjDZKvD6HKqph2UuNLNpdwA1mPMxBQFLbUKjcAhyuKHzQVz/s9MZ/pNYersZpiaGrFO52f6V
sMuP3LtV8KOworxVTurQ7El9p37JKkdJt6rjxWEg9Optw4Q9Hm+eSCCV/3KJEW2zPjTOkOQnSroU
CX2yG/2IBwfig0D8eJboRFo6Y3C0ctxnz3muNT8hp53iJHHL87+Tw6am2Z4IsHiP0kbi3qGlusCH
eiE0HwHOnGONcGi+7AcICC0sjH89R0UZJptYeJCLmAXQRcPb8uyY/pfHQUsgWspBSeebIcwufhFx
I5tGL2RsDU8NCR9Kuo2wNYIO44XBK1JAtyptwBoAGE+ISnPbx4LyayovV0TvslnzAbfz5E1cG6uf
awxeAtpMjxyWBpsV7KQ9T0xIHA/20RtTO4A0ZxGsi/4Uv/u0ve7mfmXwxnF+FLVYWvYzR+w6Tnsd
AZ2oPWGugQpRTffclZAcumxr3TeMC3JxhrbvzDFWloKwh7M+WCZxyyiLC+Xyq1hJ0iPRFtFTV5eL
dvk/T+Dpbrpf8P6mGwassMJJTTFtxOr0hzdI9lMYIRFwHUhpkURge+rImH6a6SzVkeuVlqN1LLdx
EbQIMq1rA7rk6gNETqvyCK27HpA8mTtdQeRNtMmVJxeOp+9ZUaFv6g5Q8ck441DyPQnNDAzVs8aK
IQxrbJMkSe/ROTXX8Qc0qLZ49pybSC0p4NH1oZF22h10GiYj7RKWWGPwZ+i8eLx1iNknUEnUdD2P
ol2+43L6AIZ0YBf6cf+wQuScid8qph8TVy7HtQOEwzPXAagMTB721njUCoE1IOAJGiXMzmprqGz3
FnWOx+DMcbn/DHtAbfglu0MxstVXbn4qHWUh9AN6+nfqyfm9QeelvOy81g/0cawQIne3dSLHDA5/
y/BjUv2mj9euqph63SO+fx4jZnUKzHwahcG6hZUiByLkBbfApoPqJ4tOwdKRDF9AFUveUVbfHShG
7EIhHnPTjoWSvNyPFrTv5TNG4C/72vQXbjiGGRQ3rqb32hdQbRVn8wypyhanGUXaPVqVOl64ISVo
SoTg1mm1kM1zvf+I0JIxMAGYwfAJN+JIyo4NBahI5oYsmy8mKYW332+FQIfQFyPDt2rGf8CfOm79
PXz0ObFmUJxPkB47uZWS5KZk2bD62iYRgA/ceFRwUJG/w9x6DqF+uRkb8Enxy29fI4ymsSRWUQTB
mV3vG6ubuHCLYRDg8d2yYkasQn18Vz39uBQq1v3c04gOg0mpE+TfYQeIAweI+QZ7VdAcDm9I/xJo
wNMhMnhFlcMYs+2E32fXjLd/VUx68th6Zd8Wfc6BiT+Zv8XS22UCl+ek6jLJeMkraregJ3FRb1Jb
Rety8r+T6L0xLHgqZK7DQMPmF//2qRvV8EGgGPQrAq6XnukniS/916r1rggUzU8ddCYqcc9YWbkf
e97ZZ8uazznQ1ZMy5SnyD6+IoeLmQHaPdwf+xb5SGrB+9sEnoyeJGwxw1BioBIH/V6ilWgvG4i/5
4aLJvWDxvVW8cjZBGNF/vG/WTHobucEDBFGCyLFy6kZmFzRizNvbDB4VfEKVaDyDp5HQy3bZN3xh
goUFNZRsd2gt5SrvpfsrP9RRgzFun3CYHOOd4+WNwmrdHIOqYdH2t8JSE4HXDLRkwviSSJmaYSET
CKIuQsSBeRYHeuRXKbGKFAXL+vbgjjg/jPkfbKw34oebApWkgRI3HILfCELX47CAXIPp4WwdyVpL
WULaWti6FIGGNRr0DZIVHrjcUxyQj2FnE8DE2SpOi91iNHjSMFHCKdbe+DSv9Ys8mo2zHhRPd5TX
l+3RQm/H9qv75QCDRk45ZArKC+JZQZFgVyNddgpgWRJQGKMhvA/3nhp67/4ObbYlm8wFSgdR7btK
tT3RR/ij5s8Euz23+RhOsO6s3d4xt2CjT6nst/Wfq0lTYzDj9uWspi5zCvN0xcrQ6XB06SK3mZM1
D1D0htrmmpJxYSPq2cPa3iBBtjrGMnLHQAckLLT1F+TY34OutHgMSYa9uayBQijZF075RV5b6YM3
xnXcuUlAFqHM4KOYfUSbrF/pyE9H9g34aRIOf0t0wmRUvJXjz7Ggkrx1acjxVbdnfp8bHZ+flWIT
nLfi3GmIoeeMbhfWkCFjfDNj12WJXLxW4QSdmET83ioKu4Vab9bfcOjb/SbUIB0YhOEFdtHysIl/
26pZVoW2P8YWUxD4EiP1U8Y8JEQgrho7sj1DyV30OOC/NZ6bCLq39+nBPVXXzUDXUPElXHS2UNK+
WHZ04nFkHwmKFi4s9K9SHGbY7JSPiT5CnN7qicnLTAesU77HxBHAOeQF6jEtgzH7jB1yIJEgodh0
z2PV3KE9Ddjuu8idMPNNmOYhjsGNf+TfnvY8x15m/0TGpFHtMQLpSZjJarDWgRKCKJ7Qo1A7ffoI
eFI3cFpkN/qSS0xtA7DZlYY6xSOLzPz2cnChQdYWsBXOR3palKKWMbxAg26vCrU4ID6o9ul5rIBJ
/TSOnySQ1kfZDQjok6kVBSuYANechcnlfhPdnSArySDVUU9zMQppHEXlE8yFQciYhodXGWVxH9Un
aEili2gbUj+zYAYNv/va3Tudpyr43dtTBR+T90j5VK831n/uhgxVfqzVtGlSIDxrtiTXNoAWABKp
xiaDArp/s5U21sas70DA/UbjZ1Km9sBaBa5RrDVsPqzkp7wepY6GFkoJZuuKEXIHeWDzFcgJTn6o
iptWlNhcp+kJV7BGogEQwM/7Bep3+9kBk4NCG5kTJH7nc1i/kh0TYt3pdev5zuwDYTU8eJM2rH4l
IFPv0zwyG7eiMXipfxukDax1pkYuCsnhHc98A1fSf9qGL1SgU6qFPVXiaDKE9AkDw78TGRXZdvd2
MFKxqtnYBSuqe3i/oKxITg7EUXvTZT77mZQe3w3h1RMdp+pkFQlm6hbc02neyPRW9HPLohHi86+N
mlsX/IYAqCSftwGYFyB/WMubRGgGitLSK2WBBe+/GhYYCZWTK9zWkH+dTI7HE5HED4uHfId0c+m9
9wLGuaj3EZcwh55vAJcuKm6c3BhN/d1qFDJ1aX6/JA4S201MepxOd+s/s1anCri3f5bbVKjqgjSj
75UKEEJu+WpbcW8V94pRbV4TbwznCZ8d5CHeKYwtHiHd0hqrHg9c2lihfqqICqo0+E/wj9By+dB+
xYYfzWkGbEKAw8INopytYNKq+tTKTwPb5YI0WpajUbyNYpt+tEqWRz7qrnPjfUBmtgX9n61WqGud
eicu+jm+AF1P8I3L/DJB7x4/ZUCLl5NpJbLHegeeiHilC5TRLsruJP3Ffp0PAQ7AHo4JreAbLEo1
XYlCUiTxSHtsoNlKimsgSFsau8Uk9XMo4J3Na17om9D5x+ZSYtVcSo+VOF/XxYT7FElzEcANIv33
eb6Q05uVWav1YHz4lMDHDnZtYCb5hSOY+dj6hsbKlBaujE39O4TyI1hhD2wf7N7LOB1LjAoqTu21
UHsqxpZbPDcaobbBqS5OtU7tZaZTef3Po4n42Lo1Zf9tVovFUANVBB3NOmAxTeLrRPu6Sy4moT63
Agbf6I11ch7/oB9ujnuknyNNmNNnE/NKUqVClhIK0gsWlCKGNykRqbxSVXjFJBFUjhqvzb5COj/p
BWvMQi+ylnXD/S1AzjDAVabWlnPFH+zLDWmWKF/rOWvT2O2RUBJjncES3sNmmiBvnsltvVVOGB04
jHZIcKDzFc4xvafnPeyoHKODyvdhgWPIKavgFXnIpwXqJEeS4yBX/EJiNOZKORqRddkOAeKrLOw6
l11s68nyiqxV5JcSsRSOqAyHPY5HpA0+1ltZTaHpekX4r1px7IYcAl88NEPDrHAqaCnICnjjsMCD
ldIbrlv5qgzXSfVbe5TCWc0AgjlUzRKiLxkGKsnARIVkj+VKoFlZLWmD1RZbyxVBRe7pyxZqBBhh
rN3bwqnfEnlxiLL8zxLK/9WVhtmODHqNb2bs+Gr/7Tuu56PbBCgLuC+cdWkKcQgDWpIaJXnZDdIa
uj/MubQ1Si4egclWcIXP+VXvzENqp8Z+otDoEW9UO9BgrEKWo0vSQG/bLWJA/heNkUVNzVHgAiBT
O4v/f6lW2k9jFhYOxMPG6iBpyqyS1TttuY4mMdSixNwINDy+DPJvgKohbNo18NkGDV7AYe3adMO+
ptPela8UN16HJf1xoslbEykRcknY6SpofRQMP+NxR5yOPAidh+xJ4nTYKIIJ/s9CzmCKtSZxbMbZ
24/NOUzQ/wSeHtogUbyWAu8eNkWVcdBDhSZgJxzH88Z/qnE6mZKrDMXfsdGXOEOE/Z2t5N8ywilr
Wt3aWzmpWZH6+XfEJUh1NyoXLNig5nc3+y6JkF+prwVNJTyfJL6k1J5MT1ECp+i2CkmOEOET2oY1
xSwqiILD5LaShJpwQedIgbRMocr0OjtudXJmlGILXoYaOOq7EeVDzjb5b4A/vU+cjPYJbRnxlcMF
tPf6LI2EYbtLCLVN/nlHWZSgB2h40z5YiWT7gquwYee0SgDkgEJZufOVEI6i9G7S3lI9Ua/i3pJO
Sa8NvTb4d0HWhupk/vdce5dWiSEX+bkesKPq7jgVAVxmi0z2m6BXvGiimhtiU4vbOgxGD8M9BRET
qe/dnfO8JpipMt6PF6HTosGUhNo5ucPJ9ByBENAYabzgL43/lzC99DSN1NlvjOIAumzSQVttJjQb
l4iGAXBAe0BOI6MeOyqnjzG7N0knwCjlNg4lBdiR7nd19sJMrA5evmlIMPjS3tL81T6gJjnBNs28
+LpKr4PZY4I/lT7pnQfImjAWR2sa/eE+Ty7dvjaXaSynUd6CjqGscub+gILMnZ8PVNcSsNlt1Khr
niydXsrVNGVcOKfIJR0EbQoEvlfsNncVqHfOUXWODoTfTYaghWhVVHg4JM0um92PuAvnIndQ6Mt6
YYwSigX774aG5r9dLq+hicAPkQji67o99J8f4FXSm/tkEzhPKA3sD+P7gsGTnYqJPCp0xkzJEa/m
OuxK9lms2hnPl0jjt8/hbexXaXoeh+fLveH7bvHBw79wdq5Gl2/QCinn0gqc67YQQgl+xfSAGmrZ
PXk7j566mrhp1fM6X22Or94LitQcub/zRttjuaG+B5mTT4qGN+PhIn4MH1COEerNn5VJnx/Z7F+I
pk4pQPzp5QC9uD1jkvJrqp2jrnTc5Sm/akIyskhDWIO1pZ2CpPCMpdA/74qj2sYrPSBEivtI6Zh8
jKC+SBZhOM7df6Rmr1qKwdWGJLdOZQU6I4XHYd31kooH5TU87J+XCZbCruC9f/s3rNVKqtCSyK9N
t27OY1DgGEGoVFXX4oijtTmt0lrsBb6xC3zbu++4mEjdtYSYgvuG2Gc64bxcOboumsIMkXsE+Ooc
Dq2Quzs4oaeRqjzpezx73Aepm26avhhKZ7sFe2O+SU+cPjA3CMGroRxgG/XF4ZOCv6S2i7MDb7WU
yeXMWfFMBVYnK7vQ/H9p7M7VCOmteXcRZv+PD01ChHCxZOt8u5Mw8F2vSmsi2ndJqlawwF8rKx9V
hg1jQK2353CNRAwotXAtDIXVKCOcS2zy6DWbUJvwdC4i0Kj6CDYRru16S0yILTya7Ve3oIKLe4LY
ssIhiDL5I11U1t4YrXfD1CAG5ld4zGeHhDli4hCQINSdDkfUKEVJAiA5idSmMLDknviaR/3dtKfZ
jWPUS93TS7APoUm3WwLGVXVZ8eF/UtOBesYfPGDensbZsdrCa9fj32bEF/3Ut+mE2llm1UXHNCEy
NazDe0YbKCj+inDhIbNqCAD2PznO4bM+xbhNsbytfbRdg/uk+1ZHQlxIQGi6w6G7Lu6eGyaT8c+r
yxxEgeK2EmZMU6E3kVQYg05GgiFJgcotWMK8hTdESwvcRZy7f1oVWZRut7+7pWAs5NzoLzjYbVDc
+cbERNzdap3WJzQV9vW2qoD5SZfGW3U4ewjuf9IfkJmd7epOt3vhzuJbe1fnR67dbm30IRTNea88
BpT4JPsRFnTXILOuTw/GepUrkQdpMwhb5F7BfXAYnCqpmWEecJt3OhNT5UyfyScWBmOoaIYXyDVD
yCgFXyScOArMotjIKBzIuNp0Y1NuNcXNIRDIllx/NBJk6RYokRg+YUvvkQk950Gsiu3m8N0q8jRd
ghnzYHPNsIgRXHWgHf+DEFdC42IfrGJAOSXYDh+7LSGzzvCn9tYO2WzQoOV8ieECSAchf1RiSy0o
wXmfVqkkCPLI34GTaruNssSLAWbV0Jl+mEcdJXVf2ODW/Yidp8XGAjP5n5HceNnQcHBHvP1/eJtb
kiZ3b8E4RoeZE1uWn0cmLz9cAUwjl360lTEB5gkdx7VCJVX8Uo68kw7N0bwFsFrB3MxcGNwF9Fka
VJJjG6ds6xtQ7FpqgX/gXMVHpnOC8t2n7bARoWmCKgmThLBeyNTud2SWLkYiNgYh0hrRFw7Z1pxd
tYJlkqh9RTAbX3c0b09e/3jOeXVwjsxI32ZbsKL+19f4LrW2N4gFOccioLQQEEYfS2KJ3xXa3Et+
5jkv8JaLht1MdjWaf8xOLTi63OlP2hQ799GRJOUAQ7LNfSbdF7pPKZdPf26T+Cl0K/sLKt9d+zEe
t14OaFe4NZXGsYX99e0difvqwIkuddFSOTa7sD9tNIuCPR9GpNguflAGjyuXfT8n/M2pyMQ4Agfx
rTEQjHIHU1jZ4MYqcDmkIWN3TzZ5Tl+PvQZPv6rlgHZnwm3tnmXzKs+9/QiMGgbWurMMt3pAnraz
4wmM8AYiaIn2sZXV+F/8k9xVa4Th7EVtnf7L3D+9I9V1T5fTRWBEODgBpCBmWMFG6IVSOKONv5aY
heDCm0zeswFLBUtBjix1FYbQLnD/k4IKZOuWuq7mpX3oAfcdujytfDL1wvAEP/j6A5a9EJHw1E36
kzgpDBpuj6dqVv4WiYaiasl5TF2U0eKo2cJftwUDu0Ocew/2MlPnJilUs883vBlDK0zn6C/yETtu
ZTj13WHGScAgrpIZ0oPAbWz+/YX8qZSqcAN8lrPY7ExXiJcLqMaiW70O2xAjXSSbmLgn5NRggNxb
wGEo9P1We2HvnNUpHz/WV/sSXMKLeGFMh3rg+zcMwLmJY96iI+whn10AVeWJSL7sl6v55GbKKFIY
Sa7zKSfCiV8q8dsL7Z1Lgok4wzO6oPNMauY+oZZLNji3JyMEwhf0MyK4GgIwIp13lAnFwijUgATP
cCVJqU56wmcqhkJzLhCvVmEyJ0uesibjIAYFzyEM8rP9ZfxURqNxcVVJjPfbnITcfL5WpI6AuzYh
VSfxdBpc8RQ8Ib45wbnjBsQ8acbY4aoG8YfMWQImhqhyiDoUE/oA3P6dg5zlMEZOBVF3odawuhTr
bAoJFBmLceAiW6EdWfwRVzvlFnGEPutAxKhVD6MzPME6VbxfNIYdI8ZbDfQXil63xHcTH3abIyYX
9QjvOPslVBWHmO+XGUfUeUEOtUxTxqkFts7dFMELkUo0RtEiTmrBoV45UeR/R5T6xaHgZOXpAq/d
+OHqpr3X7jua61cUEMeLmMSk/eVMX91PLvvTqpg0E62dEbDsQ/vQQ70j4IQy/pTKTCDJ8oOMz98T
0Pw4XrnuJPBtDJcaJdUdUC+KtQnPOkCzua/lTq7Cyi+j7Xeo2nvo4pTq0rj+30wKAROks7RM7z0X
FOrd0zcnhJ/xk3q65UiBB2YBRHEDgCsd7uSrzriYBD9DXbmVH1DAPrSF0ektDwcJvaXVDW1gQzjH
e9xFITosi85Fbl3ANsL3uapq9QaRzWwAQC4xmrZGMiEE4PmaVa2YEbfiOms46Bv6NI9gGpkwqQ22
ImKMJ0ldR/QMaegAhcfeGhAwinE63LbgkzGFARpDXjhkufIs82ByF0QyC4cJ04LYztsfKHVjDBcC
trcdVNFle4lexM+zY1fYuQDHWfzMmnkY2yUAuT5KwdrPgLwpuDg8jbjZS8UCOdCbv/yHXh851Cjq
Ach8in8RmjmeEnNrbVv3XsyPIpLnioyrMmSAAwZaAC9GzzTT85Bv3Fl/PLs6oMubGKkhd086MbhM
IEyOIv8ubaea2CaO5ak8Z91NOUkGMLbHlSIq1Wu7ZebXdR6iTInXl6VEbML9j+6Iovpra5poz4Dw
1u2HHA0nMKPOl+sz/vBaj6QVv6MWGT5hc9yVvZcFH9tiK1dPp2QwipCSDo9uMaPf//QPKMwJmN/g
yburClPgoIxoAotnjZ4AGioY1WH/Xr8El7ObhK3RsL2x1vX6iHiJTm2aJbP3PHgDgekEEmvtFAlN
fl4N2Pucj/2X4iOwtw6ovdR5KDSa84Yayobmh6hqMPiFQ3I7Jn95MPpSBTwsC7UPJYaCgmintmTZ
7VavAlowCKd+/D8NosCt9DWjFeiOhUqP2JRII6n06UhxGW2NfDYHv0LW81BdIrRMnDEC+xbNZ/ug
skpXda8/bE8mQx7Pt+YV/kVnoa3vGep/7hxwpauUgqHRKNs7YkSbMUj8tOEZgqZXXZ9yXAfW6imv
1xOJdXoXZDffi6Sa6ZY21asb2Ce27QDY2dcw/wVshCvgzRNaEMlEO/kXdojxUXhA9BvAvv+AVFPR
KLnYR55liy6mih9pbAmL49M0UKt1TNCuMXs634GFVjK1s0nZb/FRRaHB/mr7JVn9bHkgXJOL2T+U
Nx6+nleOAn5RzhnR/8lBe3bXvpmAi+wFieu6GArRpvCuf9hVOslKSx14e/16QI9/2u8omefrjRBx
IY2Evt4OYZ4W92HqyUBKrc+oSWnHcaHetlDgti2C1MD6zRTwynTN4YtQ0E2E8AIXdckN/LSPLFOz
lqHyYt5PDNmbmY0zqvl0TClWI8vuMEV7RtJaZRmAWRbbONz1B/t7smgx7PMddkBboIVVPb2mxd/H
Xn5uDdvni8GeGQddWItZAQm09Io2fj1+oKvMAS4TJAADPrtun8AIgl6JSSEQOfhOyM1mdnL7up3B
dfNHBwCYu5SSF1MD91iRy6D2Byrzo6xhTJCOCzzazKoPhtys4xyCVsHa0l8HH8tIYQ548hLKge4e
b8tYU2YH9iiT3pjdag3UkerMmiGSNlYyMc16Bhnet23jdSp41Cv3m4bCUtoT9yKj1UVJTCUOc9vw
bHUbwbrQAoVS6lyZrWoJ1cp3rtWKFuBE9XW0Sjx3JWYLgrrgOmQ7KtFxo644oSmS8+N/sXuoH06u
dCDeGyJDhOUuqVDP56srwTXdKV4mavljS+bvqHdsD/Dd2vSnA/nlysqBNHTtXhUpPiGRH4D9fB+u
ZDO5VmXTQNTSvuZcjnoixPCFEWUIPm50ZNYiAeBklZ5Vz4Z+fOD6vceWce+qBL+x2Oplam5zYaOz
Gu9XBZSNFjHze0rDufEAbp0cDMSBpId/gNTwtNl1GKUOb7Rg/FMgBUXmjvn9906JcnxJ7zO+/Swf
C3H0y5EuiUo+iljMr1rQB2lqbb5XrBAdxrRQG+yZycK69zk5B+Ud9sq9kn4a7Uw/d46TTmXD2WHI
hbnhbNu92gnfYdBT1/s3CRIcO8vjlTBPfZn7rH6CmE7v9zE3Knr7wNo2516Ly5jhKc7z8iphsyhT
3CyIeOREzKC7BgGBgP+hOlhY+HttMLTR1lf6xKso7g6yYJ1GIP8oUq//xLyK2a0IDnUCSFBDxUdY
OqctAJyJztKjg5AGhFf5GUAoFTCIqgvdBTpbePyIdfj3u+FOA1c8fSN7h+hDdket3dsvvlGuMpbw
jSvhHM9f6dp5qY7AqPBxt2Jq+LHMbfpg68C3CVrCumpTH+khutQloPGxA8CwjBxJxSG3WHDkZRMO
FX8grAqQMAd/QZTKSfCBIiNnjHDudGdwazkJkLn+eAtfx9y+2xnQhWcGpFoacDWSUMojF57dHQaU
bu7Q3xTSqO1f+QtDVM79Wkt2R4GKGm/821R47CJoM/pxRpl6KYyz0JB1b6oUDDmy/O7QIClD5lCS
NZ1MR5SHHdjh3Y2CyNw/D/IndS5CrX8PlHz3mCcC5KMmwJb3nh0venG4/ubESYG6/h97Qj2PmIDz
7X9BwC+CnvzBge8oHq5SoOwq9X+3ckzpM/RWLqR2NOMPFYzwyhXzdjs3btt3jO6dTc42bvVrYaCn
Jcw9eD3LK6urCj/81WRrsuW5Dl+v3bB/6QD74uvJ08sjAvPoHdh3Qd6TUrVB2CN+Y5C07E9qK8Xg
DQH/FkqOg7GTlck6kbsBhQQ00CRhj24vhvVT2rwYoyvRr+dDZHs0ln9brgMOXPTgEaHsrjsQofzv
tARrPsARyo1Ytj4rShwnkKrpDTvzAvPsRS4DFjQjFSD1SEX8+HIMyBf9r4fxS3kTLRmSIUB0Z4by
UtT5jRJEhGVqFK9VmF9g2gW0k9P+6fGj6kseCrIyEoe1n0NWiRI6o8qeTWH5MJ0XJ04+1c3XVOvT
cfq15mQt91MY4rUOd1tzcsHWReILeYaOwXdl6JITU8EoVYiOFYThl0ekFgMxdO9uDmczSpHqvb2I
VsjeI6P5n4DUXPxFXHG+GCzPgqTOCgp4rBFcvoEZ4EwFR7k0H6lqR/q9Yvr6z887s5r7WDCEQwBN
XXN7Wm+v++OvMkNCqu0yq1FP5nvzSwMw1at+GHixTF+fhfo68Kpr6NOuFaQp4eSx+7ERPcIZ4Hjy
wGyyGrZ4xPEFJn9c91PKDLVb7qhxQG8dWy7kSrdQsB91KPf7dtiK0Qj4s1K8T+xB3izln3c/S32N
+ovCq/l6kiYyPK0uQAhUHeoPNb0mJjyTmH0LDzz0B1AXw/BeXjFYL0zCgWALPXdS0WT0yBvaCv8u
OUeIjCLbEG/wQeCoFGi10gtvsBwewkru1Z1mkwj69ukBPx6IAD6fue1vB/yXabYm+Td7P6P0urVa
L598mXFP1A+pVYVHZdRgXNwNGv1fTCqAj2Wtc5Yq5FOa2zjmEzU2aYlMPwpffR/2gtNVkayG8J/a
6MDuvhZ+SlRYkIW0YlNSWwS6YswGvK4W/KsZFrXLaSAQcf4deTuKG3Q3i1ceYbm0lBnLv21qGjkq
C4nosAx68mdeGRAGLzf0Qy0JsY+VoeAEPOlyOYbMH1IoDZVpJ/pPQmcSadslYAT286dA9eosxMNd
zoQqMMT+PFJn11R3+i1lQGbfC15MMRQOUfDspwEsq0O320xZvf/tKUokkLnKo+D7XxPPCcIqgRgN
3k0vhlr/jA0NW4empPnljfOVAidLhPLPW2OQp3bZTo0DIf8gEixMPrefEr066RXj0++seeQzOqBU
MADVcjUiedW7S6oj19bWTF9Nf4D3SLCB4bsIBjko2khpcJBHWjuFmxaVehJ8ycnpnAdCpD+FyHz1
QK7uHuEcSkCbs7joIs6O18nehVhwi2CeJJ6OkqroSC4VXxaKXQHa044YL4k1L8XP5cpcVzUiigvM
ugQWHBVSoGgwK+Bu0efRs11ENUrJ6HRT0afdidyIMY3+qAC5O3eGU+7gmIay6SBm2Twwl5sqvHz+
PY1PEBwHJABW3qaRk7PX6NvreQrUOkyPpLQPUdU3C/8pX9qV68OCSL8gZhHHxIpFiLh4gNwVjvrP
cjzoHtj8jnIyUo0tZwk0DYZkloklrA4XxxmePitKcObGaQi72xeq4pdqaPYM0qROBIw2UGx0wQBs
c9WuIe8cgIt4mtvgQXCAbNpEAt9cMFvxLyvQqaeLgMr9DiPrgo7W12Tf7FoQ8bu2Z9TkX6uNvXDY
5j8nt2d0Zcwv1eJyJLwMpHEpdsAffSvMBS/OwpTxr700WlwehtMjfh+cAyIPmltDb/bsYzWkpTFn
t6wP7cGxKfNLEuShl6sUBOLpNYufDu3fNQhC0T3rJtlH7Yquc3OxkYngb6PpZPcmluKDVNw3LUE8
IndibExiea2rwXCeftdDhAJGd2+O8bDFGDtAC1PkX1NksDImL0uZFn73oWqNjQ8Iqh0P+c/w+Kr9
w2e5cftnX8aZo5ortbZmHEKR5C0ab+kzJGsCeN9M53EhybtEwUBK/6Ib+AnpF53Vx4UFnefU+V9S
DeucSA1TMqhXb1dyJcYJoKtQWj/RIAg824CSl8vnNYdXuV4ZmB88werfQpffyWHnh4Ex+252/llX
1Dhgbi6yD1LhDzkMoHW0HbT3+F261zK0KqFZrcPlC+AT51YesrRKk+LZ9XREfRQmPrK2SzNj6nMt
qMRKJxRMBs5eK3esRbK9lmAkPqUxPHpnJvgGj+77rYF1+bg72EX0yleSi7x1P1n+qCBK6oIw8lAi
ZagTke4p6a6K7KUN3Z113FPMEnRnmJD80zw5gugICzC59GhIhm0v0NgdIDgx5RLzU/lf+SsLYfGr
Jiqr4TzPqnjjbUgQeeVivMQSNQzHVDvl5bTj23kW5wg99GBsumakP8h7oXGSmOG5wHJUsa4NIH12
2FHD2+cX3H91J0CszCsGuETXPt5HOv/rTUjh4ztZX6epolSeUy5ddnxswfzKXz6REOHGV/AmT2my
7JMq0echyQ4BpfJCnP8FeVx4g0SdtVJj6LJt2IE6hblFiowbEh9sBv9xD0XPKWfqXq1Q3QTKMbIC
m6tPxZxsXomE46DwdYX8YkDy8yv9wDMSufTYQapzNsnJ4uTe0K9f9eS5QHQhMdbz4j1zuzgTtcMe
83tlJnsIw+KxHkhId1lYCfsdRk3CUgvPmKucmvSMuXRgzX4aloUGD5P4O1hZXFU1GbMtqtPT8d/r
kTEosLt3uaNxUIAhsb0CWPoEAwMBisq6C6itD1YXLFDKWptsy0WK8vPZGdmcVWNTZhW2f4lYlhl5
vlTTcFTTl+/X/8Rx3UmS+YFsKjXifzmjIrMH7vCUp9d42GIB8SvI5z7jQ9du1b0GjpqEHO/HIxbx
p5IeRGcMB/NjXR7L3+84bJIN6ctHRQqAL1UkqIZG6Jv1nte9474IIMA9F2QsGKkXDGtEjL/jg0At
wc12vAFtybghpJrbseNj6+NCoI9f6wEgF1Y0j+XPH2Ba/LhXdXbXtDmJVLt0Rvm+EpiN3RILXekX
fo9yW0FbBQrl12X6mlSILyagODiG459P02reEqVSRcuxYtp/L1tHEoKNjh/3cjZZw7lpT39HbrVF
uIjYk1Du30brzgN0z6mUCVojBxH0cJcJb5BmSeJSTKyb75YDhytgUtzpFT03Zfw4/tm2go6vpIqz
7p3LDN4CaiOdM8A1K9BG2eQN3jJIsvuJfbSs2nglzWXdmdcdnd1yqSmhc1/E2lz2cmOPuY6K+ogp
f3dHXbYHj0qVKbv1zEQYQpFu5Ui2ELLOMrVZpx67JdsgxPFVpPX/UHEUhb+AafgTf1YiATi0/Y2y
dmI3Kd77fHVMSTmdcyoXVUw5gKxwsgzK2TiTz7RbjNQClkXoLKxii02m12dhVeoVzxV4UNr38ZTf
C8w71jagXWhZTpyqIwjx09tiwTJ2BuVNqNRc9V//7oLPiJlgdNXXMvO4gfyTPtngcpiMY7rfZT5M
jpi21vBGYkuWuKRnaHBBvGjOOV7O/VDYs/zYk8XeGpoaYWhK+xYXh53gzL4vvS+0rsv1UKziBqTp
v+IgB8ap0M3napJU/eAJqslmNsONF9XQSxVFuHxfCww97uVhcv6yxMEj+zGlsnL++HAZ3f86DTUd
se56YXlxQDMhpsKxnS3fw/Mz99iTJdEq6paEZat40X8ZCBy3pSVGh59aDBU0PO7xaeK+Gslz/syp
+zKa+HldREEMDQ7SmmZOScR8EryG5BSEk4r3ZchJNo6ALwX1NPeKB0DhGZyyP2DJUGrrIn0v6uqG
UKQTpeMqiEs4eeCNDkQfs32bfb2lb6o62x+S++69dwtwnjZQ/ttXjzAjGJ37SE/EkGGdahVZbF/7
BuBSwVeIF/siM7SiAlJJ0A8JDnrcY6b3aLdsS8l5+rgkNqJdMHh+h0NJhD5LnUeHgxSlZZ7gXkyC
Lyn1mcuZk2akYhrOL6J4OBN1PXZzzTEsQOCd4vFqKVcBGUVIWFhzD4X4XrtJTRahUnaskos2iTuZ
o48PzZFbgaxaHufpkLEzYpSVGrlrfi5EgmFmiq5mFBT07bE6Gafdld63a41k45TvuTkJ/1wSvBfE
3NZMPfIL42F2Pvp0ujMWsFAdMUTToZPyepDFoC0YNIQeIFE3Pv3su4MhZ7bv3LUgi9ewSD76S5nZ
s6NVUmHSX3greJ95KEAqQ403HBSS8xd01v3vavlO766F6Of8Qhu2kt2oYXQhdy55O7hUeLsEDleT
072lxVCYSfY2G4reT/+KpN4wQJ5YN+roYJ7mBX3WBWWP65tT5Dndf3znoEuRP5ufJmVKppYAGBLg
z9cIn+orE1Rc+hwDqs/wmh3kwvYqWM7/VfHKBEGWmleGl+2MeO6CojGx1oQO0kFrR+MKOUA2+AAa
Yi38juwDKS20PdTMDNl3ikfrb7pFYo8mCIvSATEfkKLF+CSuYQ7hX1Z2xi01BAn4m+HK9lR0OkpY
kShK/EQ/r9gwN6AO2LSAjh5WPk1QszX1iKge0/tUsuQj0j6TTgU1/7oxBrU6QL5fYry8q2Xy5YS5
KelIpHC72kghOOIjEjgdQ+NycyxqBXidIJ97Wv7kbjID//rlW8IfUcK4O8DcT7g0K4xKys6P/Y9y
dVR63v+Af0rpvMIIRWgGYN9dnatQDmryxWT2ZqpxJju81b3mUps2aFUvjMeMpqDxkrvBQ2mVOOKK
tHOhiwNKqfJJqL4qoFz0c+Hn/J1zJuWPNdP3KrIklHNdyRFMIL7nT4SQd/IXv4UHk3U7XNPktY1t
6MHdOpTepg7VrITbyw7Ajg/AEFdaPFBj1D0HHz+DxxBplNOatZdNTIBX8uHjz/D1SD7p1emb92qi
PTQ8l6MMBotdvPx7JjmC8hABIAVjB+qhj+Y79tuIj29TQ60+DfbmdqS/5D01xQIzLlXoAVgGVAvr
1+ugdyoOcV8KaIC+z3id0nN+zpoBhZqv1v0/vW/PzWc8Zjuxa1+lCI9Kc/jgyomVf6YHsB9FlCX3
ugGTSIgFkCTNnHKDGSXY0xw6mTnX6s4z7dBhyhffvehGgUAqa83aWJctq8USD5FdWdag6DwdlRxa
nz1KEWsBtzDdwUpVQgvf4uu3WUJTWkweJDoBUU/JyDeeFIij/vH1z649+IypKzC/iaQVxpRr8few
yXzdFr93krba148MSAtgJgKoI3xO6BEKRnCGzCYMow+Yke+dCGa8fg384dxD1bTX9wDGwjQPcSnN
CjMCQT+CNcAiKv4TUIyQI7Dt7GXJ3kS9ChLVstOHTg0xiJSHLDcHwJlvLjgIQJrErudpxJUBkb2A
bG6YtqaMtgLjGyA+hOEfLoIC3NulR8Kbq1eFGrQRDSSQnNRbUMiyn2FV6Ko2Tp5FhaLjepav767W
j7BWdKacDoTEgUHVaTLbeduuFMiWem2MTFTDY5pJJVswE3iYrWxlubLxV2ZbvrpwicKRnUK5GXRm
1zZm+Oo9ADGLFVMH3+8RlFOXQH+YebbKw5VVm7gLUqGqLRzc+tt75PviGgWHf/FbbK8kc9SquZdO
DAXdT66WFFcG8GzmJUZOQ0tXs7jswrAHe3lqDQbU+a8hQMlMw4+YGwrKaXPGCpIYEANztbREBeeI
C3d0XW3IuTO0y8rTK7nAeyFSOIo/MkSfEbapfanc5x7XvbYFSo8/c+1wqfhCyxxoz8DOfzDit0Vg
n9bRCUMB/M8LRfWB0e7kdQV4z2Lt0k5isxHU8cjXD1gFpPqEZMRaq0pMdkLhxzou7TTVqIJ+djQe
QDfEfz/Do39tew58QgMFC8GOxJAyg/vSZOW6GxEliPcuAQQl8zP5Oq+nB7aO7HrfeWggkY2m5LB0
yhG8688OuhGhGbzqYFhdxB+Rr7tubTFLs0ohix/6I2ZXye8o3N2dfY2KinS4PSuWQUbV2RjTDdJ/
4osOjN8bWgJQbu68RwgNhea4CdXKAA7l60H+DV1xrw+BE40OKaIcxr879H8TvVm65Dne1vGa5Qb8
SRiuU2vjMROwYtGrelDHSoEnZWXkVg1QdUF6vBIo87vtE8zNJTEdKzh7CRbRog1sSRdsXx62rQOt
/9sIzP8xbuteTY4ey9r0cuTaV6KmjMb4Jsc3+5s79LnDIokH2lF88GfuCvc72WUKu2CHHfGDbpHX
+EjLJTLP3YYSfZFWjKuG32pNJmGAPWgFAuJxSK6oy2urzFeuSD9qYnNIkVrfJynXQi2h/9p4om1i
2ju1+LQJhj+8jgK3ufP1wP9Lv6TsdlFGaX30UiI3hhCtJ6k5M7WF+LqBNOKBT6TY/JYdJs7ZB6aI
D4eXGIcMeSCA10iDETAeuedCJ8qES3G38ynDn1CZnRXI50j4K9afZhEmQGMc3JQMXC6O6RGBwYyV
cinW0QMsxaeOu0qPS9e8asiq3tINYdjB1FiaOspH/uGfMTRy1LnHAfqu2L0DHl2uin1YPXqzkHHD
qdTxLK4ghyunVFu6DO6gBJR3rWImd7UxE4putjVL595VKaNES5ochLqedJFLjdHZs6EfMa13brns
bPf3UriyGG5/QXi2wyOZxKyNN35fpI2DJOLc3RnlvwaroeVknRWhP9IVWvZYe1ZVSAXDR9ACEtFE
FtEvur0X+fpmtzzEjJhPjdsCNSO7rx+9sfimH+kwueT40CovQJFtfZvMV+eL0bAC4hDGY0mndQ23
FPanQjenTWPTtG+WUvdp9ajmOYJ/5/rCPz8NvPCJpNEg8QxUNuwokLQTOFRM8GTmLS/DF9QYKVrG
MEn55uDDDP6cDVYQ7w0+UZuSvZWP3/Be4gFbYpA9s/blMeoipmt3GQPa5TXZ7BqK4S3G82kQSjqx
+vIeIe/0N+42PP6jXbBWWvkVwJ0DdEf+HyWhN7M7PpEgMD69XLCHcuYAr5Q22RrxFPwsuu4UFpIR
Eo4ttH+aMOS/ZOuQ/4OlxY7DU97Xt0qq+gwsTUBYMHzpr0JY82n7usAQLCd7alUeYG0ahD556q86
pjiKX2w0zWl6k2q3YVaQTYVymzGRKwCi3091lr4YBrA/v8x/G8MX7HbcpkZYXumMvvzHoHMASkLR
EmyLU+ZgMEvBpXGrYxRcBvneG3Tv0jQroztO6pUt1obtsblPSZU65dnHkBQJ29Om7h8pR6BsqJnx
74Pq7GZibrh7RcVt0G+soGEqSoo8Wpg2ispDrl/bTu16zXOfn8qmHrc+O2sRSgbp7VzyljfdCHvO
K/LVhz3n4ZFav3mxE+XXHdtGckM7QUxYEW21yQs8xToPYWDFkNoV5TudzhmrtdZbZK5qAiXNaalA
jXyFccLW9BDhL9hOi5vvqkxKwhAddVl2dDCFQQzuoBJkMyB0/ao5/X3GHO0r0JtI07FRB6fl/Aul
beCAi7GQiSUI+ZDIWf4FbI0VR+kAEo1cge4T8mJcc9wYq1+1FsKQjpCkFri9EvddXTYjNJi+FCs7
FeevBh2e0YmPjG5hLLpFpGwCg7UYnq9zDW76IT3XjDfeMVaaAeDiscgDlSQofxH188hOMUD2o4Ee
VCJ/BZ/kepQiDOvdTT1iH39QVAWuCT8AfTT84nqueWRaIaABUxJ78tsc7QtvT/SU69Aw4yc4ZZd2
7DWAEHc+sIrMFnpgh5ogPrCZ54bl8voC6FZZ6I55Omg/n2lUx/zQxcUq9kytIZ+yYBtDVnZf20Aw
xZnOmrQMjDqOAXcMQRM2tvOeQUoF/3Z6/NWUMJgphE15Fmycalnxc1B7r7Io0WxhoE1GbHPSzuIt
wq754xzKyCDQOcKN9d/15XaoIRMjo+mqx+eHw+C2d9JPsUqYSWAoZINCcUVOOkWfpH3cUatipCcX
1g1w9tUjNYPeHnrJcFyHpYOfL5erAh3G4SJw1ZKMR9X+pB8TE5UZe+q0X64370AyBI0YBYynDqzg
7hmL9Ou2p/vfzbQ+ZCqjIwqfvXOGE/RYuj+tRup0oJR40wVeje9vmJacXwmc5RZEjk257R4dcpoY
TY42Z+BbSVsSzvyaN3vCjFDde7kBdobAbcPFlGQ20KaiK8+uY8MZ8dqS8SOJg+nz2xNveVTGlUpq
BehcZhZ0qNPj4Tylah7+mWbJDL1+jJ8xZgKZNEru3+9Zxg7exs38gY+pTMtRtF+w4GC8fvVRGSDk
856vyBL7SnmYdz7x22GYXB0BEh3Lxr5/+B7mC+JJCJMznXVfDqEJr9mWxgmUsE6YHHMoxVoOAv4p
pFjvLRFh0Wzs6GaRXD5sfuJ6pKQCZIL0Xlcg6WM65R+GMLuZVsqGm6ggcqDSsefHo4JV+0gygMos
N6faFcP0DXXfh4fDn44XxOP42dHu507caIxoxUXBzi7eaTE71VJAE57kewAAS/y/hGUkSms2API2
qapGK0xAdR53iLGl8sfnqHpdu9+rkoi88NulGl/QhyQj2lTp5CchL/XTEW7a1veYuu+jqdexXy1E
QJnOZ5hrC4ylhkWlIvnkZO8pUnk7zNGMAkGLZ9Z9u1DSTw0hIv5mDIMdcFrgBBNFbZ7xxyykK/zA
QaMyNAlaYzUrZ82zB3qGvxTZzZvy9v8rflBeERCMVGPPJFabA/rmjdLCQCuWLqYL8xZudU2izNkS
/xUNlJChIMuXVvhZgr26djXTwDvYAhfzW7V4feq+uY0xDXQAnTD2/yG5KwNdPv+ViDyFnSI1QYRi
fazQzL21yZ70ESPqkJNjoc4807xgaXPBA7qHsPunM9vTgrXxSQw7Isw9VeGz7yTDzjxIYdMkXmmE
ij5h55Jz0jGgTmvB2tUrSgHUFaLFOIlWDRdPyObOKbs0D3aU23jW+V3uhVDGUXaKfV5GyOhD3Z42
CFyq7Pa85SgIYACtkgvP912g+61gQ7QSnFeAUcAzftzhAmYp2BeSb3QPu4Eu/M4wavex8jJk0l3f
A8ccDcO9pnTnrDtNI5Ro2Hxa31EKAS2UiVRZkP4Kq9DiWSja2G0tOWxdBCFZfR3M5HvAnNkU3FYR
wqfj2BdFYFxqPosAZ5ocT3ykKkV+nMfk8ryC+eFec1B9H+0XPlY/MUMAESIaXiPshRerKkBLwab8
hYCC/ayXPy4S7pRgp21R1zebJyHhJjar1icgBRNSNzdEGuVaWeyn6ql/12GVRZ+7IyZsKquWLaQG
xQeunQAmBiRKpUzqlmtbxwbp+BfqMI4zARIMjmcUoEMFqe/nMQnlNXKJ918fZCxRWAaoPE+eVAd9
NLXbHJvpcizOi3jUIcITWVbmV2OcMB4RhQRxtMe3iI3/L+YPfC/L9W9xRHjTYmTIZQpVIgxQafNl
6JFA1/dAhPYeC1ZcOiM3KIxIM1p0zMjIvtriMas23B129vb3bN2RnPyv2kcPkmAulPW3erFX/zMJ
Us+S1dk7JPeOuJ0rUsToKFrs+hQnC4B94AIOboVBH60GhLuIldww/zMfl+0ZPBbbdN/zIBcRC+4P
0c8EP6dPbJZYzs9Tu9EA8xTCcnlfqKXdfm8Om0oDkcKhb/kqh3D7g5ZK6cgl9tY6HcHvcHZ54MQ5
fUkGNqaS/J0qpTkszn7+2cPP9l3GR27BtCTb9J9p6GHIM7seoL/RH7E+ZHYP+tUwiy1m22RrPTxb
zmk50FwOQLSeY2k0DEpP0tu1Uh6YYXFkwYHIIjCytBy+4Ukv129rSscohmsRvBPjx4pvIKP0Naq3
7CvVeXzDE+lcFi3R1+GlduUk7DaOOwivhieUBRmdRfGzPx2uOmdbOjJmSYHb62UCjHllfcM1VDBG
zgTZ9KbaOwm6HsqV7UN1gUIHEYEpJ7o7RSTf0NsqHOhCpKgWFYKWB9Mph67gQBM8OGrsLd84g7hj
O2FTlOso7tPnvUAZIbhE0K5YoBTjq5xzomTPEh4QNHmWbKoauDbbdcupOS1LMa5hF1CyjLZiPA12
tDhZKdUhW8APR5E4u/PyKPTnbc2gWpVRVBzTV03SBEClLcv+3/VLUjl4Wxz+rHg/PD+SduEvITo1
0nwxpH8g81D9i8SibSCRijO68TUpSEtxup91wpAnMU6Gm4akAIgkXgxSgse/BXqqap7XNbUT4mog
8/cbH+Q0C4FAG7xr2fyFDi0bXQ8fjv5IxSUBHxGJlmCtoUDeXD/B5w9Arkn1qDKEQNJdslA6krdG
ME1IYmfEXtMWLWJ0xBjz5O28dzG28e6h5chk08qqGl8Fi2QtKrMfRb2Rgi7fEFqumbBtLvTPpGKL
1vy/xhiaCezLoYDq/NLqoUnhEzujQkRZQiuca04YrvOJaO54Za7Gg4fNIFh69h+OeVV1EnWALDQk
pJoYyQp6Kli0Z0ytIfAnWrjwaF5bRVUt4Um/0ogERX0z0KvWzQdiDgmmP2TEH78Ec+P2mHTZ4Y1C
3uBxPwemsA4TYogmseZv4Q2cTXouF4xCaLB8EIf+883A21CQ1Pb7ZfLUGdSpiUtSFBQzGCc0bY3R
8+828YdKfSypNZZ66nSSfw5QrJ9zFqZFu2wYrSEJ+BA0oQ51ucbCoMRcmbAfBJ/Sr1h2MN9c1KEz
HRptnpQhS0DZ6p7KDPo4w/rrfO75zHVuY3wqygL1jD7sojOQCPDZhkFgBrgVuZeImkrpNZzkMGMn
gg9v2JOXih9hdwwEJIN9BkhlEWC7uNqtZ2jtfTtQ0TpH/yv5/rVP1Nb2u3L1fJQuQ+XSwNDCf/gv
0HxTob/QKeK6qii8MJAtVBCAkmXu6UETL4MCkAJLmn3mw2veFG2wMbRXEibj/uTYmM0VRgPsuctO
Se1VQKkn4pzsN2W2U12y7LbFyT3jvDsTF/soE8u3XQobwXg1ummvMWQsUg2NaKhSP/+1p7YFBYZ6
1bq1LGeXiljWxvrSAr3gHmFM9pToeYUxYzzYFEmG0aIczbLiiH73z8+bwGwwup1tabzvj2rQz0NV
50d5bfQDW/IyTtsohy3vfB9B1wKX1iLjLN/OmTEqMUeE55eIsPH63nIK30XAGfXnytoRvmSTNUrv
8+CD/SvDpgn5oriNsEOXiNW11jnxPvSmK6W7eL3uh1etni/6sO66cJSuWfkF7Yt+ogwNhcEd6yzg
F8wu48KYCE7pgLnr9MysS9Sgvwocixr9Y/Xm82oKtBQs9Gd0cYXOF/bGvTOro9jTJ3IhIfGmaeQO
R5YqQ7UWLUMc/Gc1ZmDtLuJkmyDUsygC+LHhxNm9DZ83zFEbdbzxIufzOGuCSFev2DvTyXvu+68f
kBXU9xt6LCF1PS/zqy+B+pSuSexYjKIcpUNxu9YLerOnWYEj6qjDQ/S6agbeTzxZzZuivJEA+a9t
Kzsg0goHqwjrhGheBS2VmHgETlx5t/DmHXvQ1ZKG48p1nAy6VCjENAtADUR2PS4yGS3bMaDuUTBL
IFi9Pobaem8dK0BO94sewJ3YntlwFk3pwuPS9HZ5GuLidRKdigsXYMzc2WJG/OLtMRa7X7md5KZk
oVuIJyQae9K3U5it5dZkXLr3FpBrzqD5NFUTa3bEHBsXk6A7wrI1rg+Ew9GFe2B6AXxpLxdtudnk
AZbHL+VGFI7qM7j4jXyeFs7JkGM+elgGl96euXN/54IshCjMd1568dtCWIJPDvThdzRzox6kM9v3
44E+fLvDB9QFLT+byAct23bkbpPzTvSIAzyamvFGJbTqlqcT2bQcmMdeG1gIuwOj265wWFu4O2e7
b8/X3ROLtOulbge3zg4zEpGci8+lhdbTAshENdDPPvgt0VOrdmk23UsYkYqHDwm3AQPtIIeFr8OR
QQV7PoUVbn1G1bZH2BjVkuukOU+uJn7i1c29WmO9/bRCuuv/MnBsPJTFgASfp7iPruLsRBfxTpgv
jswKdRPDiCWHThEjaItIpNgTM2xERn3HQ5pw+WRS4OtPkFj1IVtXIZQNqT5pSTuWrbC3OMarmaxI
/LePcM1/mVH5K03h2q03BG1V2/q3Hx7Yw54RLH5kzgDaznRa64OW+ztes70stMbzvXOM4TUzETV5
x584m4AMs0tnZxmBcTbMWo2MupLM+/tuVWusFYEGXnEW3R7hl896zKVIbjK4ZfqNEtNzEUK6nJeM
08fbg/XbvHObNLAah3n3TE3VgswB+U7l8+gj9uGKdFZiOYwASrd27cBwR0WwJzc0RpKsqc7pdj/i
L2AAwG8EmAhJwY65bPzhhvZgAViuUu78jzpN5kbSZ91f8pCdunm4psAposWSVX7g8G1WM+p0AMf0
9Z3m3XAk4ON7/4+43scspwuOqjWHB89Lo1Q9RWJqnsaoE/Dpjlffo4nEsAcciedVkaoOGWwl+4QM
+XbtVnY6fDN+mUW1dZu90E2mhWjUMyLGdVIrUyuA9GqJxiX7h7mp6vpzHJHgLv0KbOgB5UiwKX/y
X9aZYmk4wbbw96YtDT668TLjYwlTqeLcGNeTOQlNuOnMKmooc2ImkyIZp/I1K6DgPLrN48XCSqmn
pFBFVOPDNRUGEE8ucUU/yLHOt7gJMBYqGl8OJh5QUDR27y0g7k3UjodmGILYXxUBnZk3+MKuiGOO
z/DfFphelMGLufUw6O3PvFrEYuj7KIBVEmOqjZDyUAvxBKlJyYKZ5mj/yVPQuobLW6XwQDnt3v21
XteKlbxAoq/cjNDr9QYheGBI27CF9jn7T5HMg9advN7m5pBU3CPVqHeLvPRpAJQTcR/3wamCr8hd
589bcKLNLcRpEj7yNh6tben8U9X7uVTMYsS8qszvCLdNhH1BvTx5/lAIHhyKwb4phdpIECAmUWEU
yJ0MGfPS8wtemSsx+gd1JzDZTOeuBUZijhMjOHOwgVRkWFzEHOISYLKDYQV0j4mvRRQFrdePo9r2
b8xrNnmd/StzhvrOfroxoA9abhAcmSYczCtShwGX4wjNT9GWyOfeQYkNyKYkzQLtmhD3SERNm6oU
juH5xXWWuAg6cpyIoD3GAkF2IeMrVJHjeYUHr9jcickgbR9dwbXVPRN+ZfqHhCEupKP6auSHh7OG
VJYMeR65X/0RNk+E2G22jnHeEOL3lobv11UObzEhTcvJ7B5C8BqvT362WifUNtln9gvISwn+lc3S
7abveSjonbVQAuIui2S3eE/LvOCYxeFgo+lXpEM5W87TLKQ3TCPVrJTFzWIw3T29ntYO+uD/7T4W
5ZvtNE2kmQwQnqsVF/LdYXoXOrnkCw6rp6FKXxh1QPbSaE1ryStVqkVmt56xF3SGOCxEpzErp1EY
ASlUM1f4QN/XGXzuza7Ruj561MhQ4dubupl8Im03aUEbcZGLataM/Z2BC6Gf2jQjxQqynP52i3/L
CgrMkx76ruJgbjozDgGnVKDEXsjlnFSszIZOTOE2KXYuSNvgfcl0GZWxqEYRepJggm5ENuryGAMi
cMk+cu922m+meBILHNpJL29RV2jZLLfXbBVAe7fhBjoNvUo+afVDBK4VMzBoG5/92lmtXSaqCiDH
vFv62kRkFXxUYy7al7hmOo9IiIBrAXOJnl1sKirrWg3KPyvRE6/FuJeRtVsjBragUCwMvqvB+0Ja
/6ryrPNJE8qBHz3e2SexLTRe2Bog5Kv/vc1BWGhfbhA15OqxUqhHpwJf/g3kbavokmVuV8Vth1Zw
WsD0gMjN44LP1ekgglxj2CytJ/lQ6XlideBef/mP39C/zLUDNxabFx+jmEFijiW5xI/N0gs44lbn
Pd2uVcJtUM+ZlEhX2yi2BXdEMz5fS5Lj84djwCc/L/Lb+AvSQN5HVXlYjZSbCYo4o60uI15fNtxz
GL/2EzP7eGn9pqeun1R7bschdTjzgVQ+W/HfJAnOGHZocAZf+F0VCWDNadPtkZlI7Pg/yH/0gqiE
ulcIkp47xJ89GAyS+OGQgq1i+zvePju0hVQ3Dgkwz48jCRBut8KxchxRT5+OG34CuTS+UkoAb5v3
J6m79XdQo8UBW1VFblacIinB8lGYkf33m3MKmcs5MPAGn6Xt2gc8HXD08PfDgQQ9qS02gEDuSUj4
JHCTJo2Qz3I7S03K0aPMte21R9mIiWwK55qeRrC0dLH4PERcic8H1hPdjvMG8alfJxxpg1aTOSut
ptRzQamj5iEu4K2F7TdsOSXmuZxuWSr+TM+Ww2+XjBr9AcOG9zTFF/f5NIjgE+aL4yYt1mUYYurf
r2c0sYAsNJfkD1tyEFJ23FA5lwaYgLr4g5AnS07DjYtw9EJGKM+Gg+LkyBbRIUXIAkZmLos2E2py
HKuwsfBDvE79Fa4JGOXmEZwb6/kttoqevdInKVFS0WcCk2/Skt5Aac5F461fOxVgGGo1O8Zi1OxI
85AGaAV09kkqN4VPiImLss0I0ru7jI6r4dGXy4k+0VyT3suc3zWYs5etQ6B7Zj0ceEbaAdepM91X
1EmdB65hwNvQDmeooPTZIen95klKRrEJ1xIYRauQ2uY/Lq9F4JDDWUNba1Q2iP2TSv+HaJoQdsC8
9u55iYZTMfUr7SJemCBnC0/8mVieu8g++j7Dtg7f3ySjiMGICsGvmtwEbetHyIrAICCPanNr1jVe
gj3CmfAjM924NRdUxdH6W7aWlxSyJ8GmuqV2hpKtk6iQlog7NjVVxrDPHlWKQDbQbNNcdTiJMIRy
0CMWmYGpg50XUj37BhmxFxUmP+WgekvBdwfPbY6qNFHf4l6luXhtfhHe7P8J3PNXRbzI5CWCEUv7
fpSqG/gBrIq9JNqYnWTWUqBfFHLbBxx4OzbW/7MRxhmCwtrDI+s61MnAdBfklE05aFihmQdlCT9c
vQPfi+Nevtsz0BzOHZCIaJ5fc9qtS9tpaxr0aDuYC4r7ZxbvEdUS5RwNRcRhZz+FVjFgZt2c1TVb
rzBa+Afaofh6wdoxRh3NSk2wQHQkKgKz9nJHeq1eHC31NhBnS56OkwlUlOWtZfk9Bc0oVtxtDggd
cwtqkboxxgJHJcnOSm9GqlspmXdtSr1wn/Dzo4QlBdr6NCRR4/sAgw6utyD+LgvqHl9+IPGvcBMv
GnmBe1rcW12W3onMBEDHnZ98Y5L3KA2z/Ndgavz8Q9jI+XK/bdH/62uoonCduEjGm0Ab6FCLSWuJ
8llfvZlxOm3gTrfrkmbjudNbkHmt0NBZC13tCJivCwBuuDPiSwhyMNIspnPpuxnHWpuH6zfT+K90
iwRWvuBUKFSlh752jLfdOqS8/PXCcm2/WftrZIzDGcGLmRRn5Wsz0OvCIA1ZdUh2u6yIWnLIg/vx
o19R22/BTP+egPzzyiLHm8XRhOtfFfK69fMKVgcfbzhFcH/q8WRTj3nclmwtDGyZ76h547Dyp2FQ
uIhP93nYmquYCG9vxHkqNbeMEdTAm8eGSweP5J3u2SM+9P0/HLuTpM8VbB0GSHvxqwClqiPw96ZS
mhdhwgiKKvZz6A/3Q5b1W1DRk9aGcgTzrwaKt5dVaLvNU7Iz6hxi5wIlWQ9fMVcNMpVFzB+KVbSR
tBZXCfsybQ+2m7E4p2W+D90TW0usMVv3wJpJ48XLLJ0Rg2I8pZzF4S/DwtvCiVUfYd5cVPPmirij
eL5+z5Ip7xjWzl6B4R0Q5ue/QHGY4/f5SSSJFYlG9J87oC0ngy/1TnHi0AXiovJayZEvGT/86bfU
yp0bfmqY02sYU56bkxzKjTRVelsSkbTvKFDVthJ0/RMo5Tfs7cjpjZeeUAq1JUjAUhZ2FqtCf46B
jHxHiO+SeMNw6C6C6TCjp84uoMSOJOBapTTIa5S/gwBTpd0IWtkesQATxjsrNs3ftUbtAKkllSUt
415aR2ooP/ryYs8krI99E9PzFdlYvr7owZivSKVHuTbwkWpsHhWV6hLBbBD40PP500leooTM+nif
a7FVrkccBQNXKr/53Dadc23U00t1wPPXOB4jKdR1cM9YhEzeibKPlVz2ojMrJM4Ox01+I5oUMouy
ZCXdceuBWsGwk0wXAp64dSJLlQWqO4FBNMNJ+HxEFVSqDCrlxUlWEWpdGPvh/bLdjn2WbkiFmS2U
lVqCpzoDDVQpAktNR4REn0sTaq10F1MIj55Ht6BAV9PKyf6GKOzfbqeq2n42hb6/iTwVxP6l+sVJ
if9kbD3P0NuPcpdMH7MGzXdyHWg4kyHAYQJjjeNZnwDTOFDsRMAlsg7VGAT+Cz/j1YEgl+XItnoG
4gGRqMrriyc9Doag7Mhz7zyKEosxEPvGCsIg2uaA1Ht4R00n6FobFXQk86yAzD3AJ3QyKNeOrGZL
RXKsD2s/aZIodJyLAvC7s4Tfq7o92/3xf3dNFwDPQa2xWGZXx3fAkVMXyp8qTkW5vHO3MT1dEQoV
YQyrDQujY1lYU+iqRuHFkPUBAHycZd6xBmNg/EUH693XjNlXVaZlcVPfWT4mR39Zcc9XjjQqof0s
el5VCm5534d4MvvWGmiEO+/a/sCH7+Km7NBBesIhPRjsQBQHTy5elVhSXlyW9o8WxgILflL64CkA
GxfamXk69WvKrllFujl2TC1qGvzzNS1ubgvs/pLoFyebv/iMfveK6dGYSsC3vDJ24MTr2Lm98pWs
9M3MOSyqJrUZ25WJSvAi4tZUgjhNt7e/4g07bQ9JsntIKf7pPq73Tk45LaU64geHTigBAV40puyw
VMF6K7ar2XQbTCjUyl4OGyn+9dsMnJNizfXzRrmKye8hmEn9vSVy2HDa9Ky9fqvs0jCo6UsVetnO
rTYCBYWrbhIpdKD5Lt8V4RJTdUqRqcUXzWlFo1me8mKQ3DdsnWCpUo7ACdYGFpRsqtvVcs3SU6aJ
l+i7wZFyHYYcxce7B5K09sxoYLtb4aK/PI5Ps/ZKcz/jbABr9kKW3rvrLdss7QnIijLm1sydi7VZ
KfD3wCtc0FQwznc4LhLsfoljRS7bH5J9LodulNtevetOILNXCmDtXyIaMR+gM01wkYaKRlgGqwBu
D6CxCNBlpmo9gd63GYAEunUHtvg4akkcOoIOyIGh4tuWtATcc/8ALn/2kBOpj/n6EwK1rRyrESUl
mVfvlE93nDYBF9nCxmz+rMiJPixnJ7LBRRlUV0AVTCO3tzykn1YGn3ghQKk52Z1vceGkL29aSVcK
PlOP2V25RSfLCMVgNQ9+IDt/VpaT5mmp4dxqVy57ZKao06n9kwbdgRpXllVNEEerHZeLbiolf9fZ
VJNxb8c4gEGNMOQPRiLuMUIdT5CHm09chHxvpqfCV5LLKDAuLChDptWZgstXAiE3vacedmCs38+M
fqiTTFIuqNYmY6vM4uaZb+0B8zkxbZhsHbWS3/SFF8D7TUxzlxe9NzMLybfLkkDKWSaEvFEMBQ1F
kGb6Znb5T997WwAMlUd2sQn5+CMFoDKvDWxRGYiqpAihgRr7zBdludzBJL3X1/Vd+yfZEl9QBM7G
RGep/LZSB4Rqf9+aquv9w/2mbBFqkhzogg0R/l8GJLlNu07esdNPKY41DSbyV4LijaPWzDiFkpBl
WuBlbLExStrrvmyBX4xY0NSxpJVMjn5NiU8WOoNho+498v85qnjrWRrHbJ/IHIfzhqQl5q9yWTUX
Rmj5gM5YB57mpCnGgxF0XdqnoAYnvVFugl+gahpL9Nr6pQr3a5clyPQMu7c7rVG8t2CumSa0Lpmr
ci116SHpB+k1BrqcqzedfaoUuxfXYbJMjiFUJT+2eHCRyAELFMYF6s8wtfLb+la2Aa/osfyD/P6Y
q+vKI80M0fJYnmtsw16MgFgt9hpupyC1GnvQx94yeI5OoagKDVyZuryYKRM0eIpPqhoDtb4uq7Qy
QZNnSQzTFC3OuPuVGUHoOQ9Q2qbzm6pLauuj3L9z5ZnAzPauw3loIkyddRbkDvyCrDN6Uk+w+Urh
gdJFPYB3w1S/4UrO41RWPDnPRi69AeGTaQ+HtxJwE0UBhfIzYFxnNmOz8qGmhppFXP/wVYXgbV/R
ArAuVeox+QJ/UAa6cdvGYadey6lHC3Te7TWdgU28nDCrLeNaEMtjXhponjs8+5QP1mQggZL0p1eR
+b5UROYI5aXnkvbNE2iSAdMybsg9E0iVgem9D4WnwgQlpQzWWciI1Pdq3rkXVIh6vnjKStYPDOiR
c8joX5GiONkvy6ESBFSlq1/RdeTowYgijclEfYHrOMvq6m7+yGXMEcBBUdqFW5fcL3VlDdvo2cie
fwJOo82hWPBQD5b2CVM8PbmsMILAPSElpRZVCFl/nq3rKmoLrlKvNt89TC6CzI1xfH/fJMNvS7NR
hbyFibyNM48MoUiuqcLe1kCtHC9O5J4L4h5uRly4suofPwyGW9GerbJhttdXfRmwAuvZDFqKW2az
WNDFiS7WrFbKp8GjfJaBjLOMpTFbwOMkhpbqkwR5bZat5bhKdHPPcdx9Avr9rgr6gbO1j+4UZA4X
Dii/eFUJrsXOnZ4bvZYtO/vPaUcz+DtLEviJOHPU+rGa8XcRDH70a8sIKQ9ek4WDPnavWB9WUnwG
sD5SJUuFqxwV/PCyAavAhtYwbEnjlHPnMJK6IDgV5hgiLtGupZ6DbdYU8QxoRjyWxeMn/xvxv4C4
i8NN+LB7QqmS9MfH21pYOuA+XiOwZN47r1XqcsN6jRDBaUjZrHzcShLnwaH9hERzPt7rGYhvjpb5
8T5ExFuG65gTfjrlPuU2qcUrihmm27kFsTpUIPN3x5dAg9SLUiSvucqclgTlu9F5B/dtH6JwhzaX
usUpboqjdraJr4/czQjqeAfNrqgzMzevTVWHSbXj62S7tMormqPfVkhTsIPe7uOYpqe9JwPJ514i
QvEZQs0pNpzPHC6pNOn7sx4XmEAKairclTvfs7rEfmmsy6W/wr7shF5J4dZ3n/ubUSGqFqsjUc8L
sXWigTOCFh3rUpAJWvJAvtDadIj68V7EH53OxFJXLvCF4GefFKX5ysEpDMunShYaVPXpY2Flw6h/
T80CU0Ryg9jt7TKqIID5tXzafUvUl1LyoOxbXzG/Ye7MWPk6kEXwUm8o68CDjo0eGJxrbg+9r+YC
Fh/rN5pRsjMmi5h838Pj1iJyWCZims1dIBnEP+58JifPHJzf8x5qq5rcygljaw1LUfDCIrxx2jJ/
bVDipqOO8RlPHQU3zhhDiVtwtLPeZdHWNbY7dedvxoVMJBtVfykyIlXsdfsp1fn71lLRqPfcC5Sw
kF3GI5GkzOACJaAIIiLPHaeVO+brEn9GVmZCryCCeLnc93EMjcZd+6C17rc4PCbXZgozp5gJJT4I
dSHg+6Z9hbuoKLkjrt9JlVFo7rqHGXQ1uiuHP6eQZe9P00HLb9lL08CVWoHR9AFotvNCst6ZZ9PG
U/ClbGPXhwYFTuGxrhuvsHxHLYagaRpsYxGfRb8TZwaJLUMaW+o71djHlG15pTRLsXSS2Yr/560Y
GQA5/a+OzmQqToyojx4N0SPbHUrPLOQJqE3hYVmGhbZrmk6OTuvYUcL604nb9UFWbPjnjlxRPJfZ
coptFPOQiMYaoCAbc3GsT4eY5SR9SghsOInrMkL1B8UyzO82raFwgvTI78mL+lrd52nreIh6aQzE
kPej7QLpvG8ua7ksTFEfdFVhoPdIXAsCkq/+17ZBKBRbNHvsSzy7G+taV9Vr6bQ4Q5pFNyqV+hKG
+PNyQvkoLPvzhQMJxWdHz9MWofgsQusLYna73DI0gfmUddmh+L6Aswj/+OXzZM4VSybr7yTQRjYV
a5ptS5io7Mv0OIYY94Kfd2gG4XQMaS7m3R6l3ZSrDIDn3xn6NnBjEMCmg9dxV2ppoc34GicG10Bg
VxVRkCMcRXlKyzfCWqLYLcW+heKtm7M2XnCQQsb7PhGsllee7R7eWTeh5ODar9Ots90J1iT6bS+z
Pf8Vo9SyycQoZSQbSKnOZ4Pj6V7YiamhsH+dz7LuGdxKeJ00LV7kjlM17S2YWPZ2l4EWKr9WQO3z
Xo6qREHpEQBIRktw1K5RlL+wFyp1aICgq6yQ5vQQmm+U7hCZrF7LcWWpD4hMIOLfOf2NTS2ExjQq
uE6TVKuMJF0aBBfDsixCwFZKGKz0aOF6A+CSZnvTLz0FnWFWIojbspQHsqlkCx3AbyxRd9VA4SHd
kihySaDleLvP3R3tU0KTCtyHk9BISwl9bXMOKmlwEBYC8a9mpTD8xrKt5UIDc4EwnD1p8caTk1gE
YH1JfS3LHKAdOGaJ4YKdCZf+o6DzTOL7J1uex19OAvqjaOyz2EvlyHzkxsULrE074c2svywGGp6w
H2GG7h7O5/ObG+lck4pj9YwHsEme4jHmKwt305JnmMmdk6EbATc4Htcz1UkqFilyr1pQqCtbsTG+
/6y/UlYC8v6+pGZpMWNzv8S7K++6hCwLY+PzWVskHMENQ0wP1DKSTPmIr3y0NXopb9cWeXtIy/5u
AiOKseb9QhwUxUv8jxQ/bIu8/Ssl8l7qYog5eq4Bp14auT0W3/bhMzKUt7T7qXNc0AH/Oy2bUKQ7
5P5GfUaTioVOie5Li3pkyeF127v6T9tIdcWN1S+15qV5Uqht55yvNZCXV9nreyCjwwwGdunSSzs9
t40TvWDZh0zVjpkTiWmQQRQ+up91EU7aQYiqhMXTzOb2G0sueEnA5idEo2Y3eBimswkGwpSrANNz
39CKJLaY6ieIZu97VW88ks+gzn1UGukQRU0Q0yphN2DC7ICV34YMdp1BGaR/yfpGCjA6R2vwyGdU
H6n4hfVYZxIfffpVP08eTGojiIKHMaIF/dNuuDbDSc2TrsSSIA2L6VkVD9yYHMQxJd9o2y6bxnVY
FGsQP6djtmAr8By1GJwYa58XPMxxwef7oJw/DBuNNOplZ+5ZrlLbsj9GQsFPIXsqbCCGmZYcsper
/FQ2kEOLnTpku+J/L1Iq3nOKP3BjSOxMgefN5OjnlrLTrdz3vIOmwjFguvKKLsWRYtkdVSCPrheU
l+8wBDa32z8tFdhSrxC0hWa/SE4pgpyeTBbqWTTphKs/CQ3b4mpI7nn7vY44yo9fVmGlWyJKkk1P
wvUPVbkJEfcbI28JaqVNilvKXsR85WKdwrwmi4jp0Jp3KQmleOXACFsy1QXJQ3rBuK+NN/9ZQl4W
dxrpuY2EPPio7fbMfd/F8iTr40txJXsbbf60EH4McXFx7P89V2ZCSqFsIqr6ZgamMPQz3lAn9o92
aIZAVHJBjObnNL2jq8YXFi9akigB5c7qw43uTF/ltJSAeFz5CIJ++TUp8spooY+U7DLlUP/h1dJM
Mm0W0S+pR96JL76T2Y8TKzdfRkEyNxEP85Ykwn17J2rsTCBpoXayhnWFmSlIUL6o2JkNZJ7ex9FC
mwX4kpPrlmNASRV+54ZWkUBI5Nf1VCK6U7xqqkh2JV3kWbalj0QegSE7b2L/0QNQtRgJblm4lgDZ
PQCLsfVrKsTjtb97bzhr01RHihvayQXraJgQzQ2vEuW1EkpcrVQ2fepfWU5CwpiJJloaKk6G3NoV
SLTdoGFBAjpCEupHfQojxGoreVfKTSlSXMi1cpfBkn1iOcrGDtGVVA3GoB2dczdzft13JrPvzmwv
D1nBP7jXpp26UaYu5Tw/w4tGqtGICN72WE0futPNtM/K6jb9RQJx0POWOuUw5mJ+gcBb7pf3OA3D
KsHwCvgJ7lSP3yQwhP+oRcV9yiR+E7Ip4gGaHnUt2PircrLKBPqGO+Q3dvrj5ba9xT8mrxWP4aco
ItkrdIGAYhLwiBxsalU9pPMRLikR/oarC1kAYVHraNZlIa/fXPmOOsFQSG6xbFMshxy0NNuTV4z/
jDQWwaB+4V6jobs3mqte6jDyw8gvi3HLt+tCrS8CHehFOs4HNkyt8dJNXI7Plhw59EvuTkhHsbZc
oZkJH0G+WF4kI1uRCx8UOxXF2jPwooPnYF8QbQTSOnQIzBd82kBcixtJwVGaZWKkz/lWfVKmsg4L
cpebBLzj4Swv6Ji0nWdm91ODNFG3nM8CCF9Cv6QyihQMmeq603369PJN2JhiRGYO8vtymO5bIGzY
NJmGpOnWjnU1lpGkgL4UIY3f1c9TzvlwivPxZnGcrmohV3wcnxw7z5CjRtyE74De8UNcYE9FW5P6
Fv+YQLxRKbRgdPvjdxJ1Px7vb8+v4MKPz+X+ur0y9DQTTZhb2lrEsVPBSvXJwq3OZVg9AB9e0Qqr
e3zBELpcz5O5TNjt1CTtRNbBV1KHO0hwT6bJble4cZl+DYKdR8CE3fnoLlAhnzrF6MnBYkB86v8h
kdkHheO21IlmJr848rY8E/6RLUC/NAJJnI6DZrMd8erZPKnVuOrb+g77qL7r8TSwzWzB1X3uSbdG
Vt9IKuA7K+zgrAhBnsvcFYBPA65fkLnmjlK5lkwJX4WYY2EfUPnPGh6xnlhGgzxHRqZ9cO9QOSmQ
kKsSBNunlXJgPAW84HmhkC6x2+miVjjfUC0DKtALutTxBLEz0++1kvPopRuzl0HNYSURsSzL5dvR
tqBTY4h4geQHDyFpD7zQfRpADI93IiY8zroTuGUo++u+sPsGzRWTtDVSHMDI/XJeL6gy5kGp3aR5
9tnJBKWDz15UbdmTceMI44FmpMzHKY8xy54QhCPThIY9OtxMLpHhPcHv4eIVUM0EXKqNlWN1Qp83
0hDniz+TjLjon6U/SYlRXiOw+npmb1W7qlH8sIQp3S9FG+7iFS+f4JIOFVJleIyZuXZIw6t+JE2Z
vVndey6A2FrhBqrAsU/SUlZaxB7TGyqKgIUhRIEFdKdHate6HFhQha9nngseLe6YhdSuOM89FFob
6vwB4LSjCRG7HQW4zN9IyAJVlgcJgOvTIoidcTKUFsHs3NxmbcHLc/ZAXttVgqOf0OxIE+1Alexn
8ejWUYFQnylsv3rlsisFTglVC0RwZi+J4NsyIjeWa2h1qCkINCpc4n0YyaVBO74JK1fbBy6Ubkp+
wJjKdtEcay+CCMPZaosig7JO1XsLvXVV0RpDHbhXx9vl3pDBBMzZ0qw40aim7aknt0cvibF8QelO
H/7a1rrHMYdk6XIfAHPXXvjWttyoiNzmJWQFSHCrm9GDNH5aFFULx4wSjzOoIQx5rTn5p5gBmn9Y
I14sjkYmemMPxQ5qCdR1saB3ui+eL5rcaiNapONY1aGfZhNpjoZcPtYBTy1s7wl/e0047lLN1OYz
F1xw1H8Dl0324VUDnZE3knjQFc8T/jKRazSwWDwkQ+t8vamb+qRDaKK5CDRBQkZf9fFLl7RO8Cts
cJ//LEh5jilG/+kBpo8utBuYWNb0Eey6rKPZaJckry9yEeoBhlQBwBVXd6Yo4FdgAfzhq8y5Vuso
bVeRqimvE/cDWnJidgEQX89xr6GJUU6PifcOAj/FrhSewjxhN06I4VE2q3FPldlLTehFt9xQTfzN
kb981N97xE0PYgRr1ds2s5LJ01xfFlORQXhSQ92ywXihklZedyqY+WwHbSj7tKHDtIQqQHRBFl1B
WQmqyluomdaA6hl5ONc4Srsgre/afsOGVGDJwDcZIiZSxVRcXpQqThpS6sd9aEeObBn9XZPEw3s0
UzIDCNTeOCkPoR3xh/1m5Oxd3XuLNEm+x8acfJFHd136BzrAeYKQnPFzIcKByz4LmAtm7ColaPRS
T6yP/cE5be+4Sht5JOV8j4L9+2okMIcXdfEeu51aSXkFKdYzjbXLGYAGok4xAYjNSByTjNz1zeb9
/jzo13HJ6kOs8XodctOuNNmIpLFngUetw0QGKEhE3sBKYv4x77JM6tHVaj2VlOQWgwuzDutWkwNI
lWyrcZebCwN40EhJ5iqmDnTITnjeAGCd1fTHeObupAy5mHUe4sn1NPWixYjIDYBxSQSu8bTaGjDN
kN/us4YJPxxUT8vr1XYk528nCR7Vb+9q54cfTXnWNXlrzkEQLZBKNVm27fXYfdP0nKB2P53OaS6/
ZZmKv6n8sy/9QfcL0FgaTVkR5NKlsxh8UoEWAEiFdTW8+5psJzeZFET1SakfXTesYQdFgDMF1A62
sSputc5UAYJeiiRyRnl6jUlA1BTmRZIn6d0zXxdK6+/cup0yLN/1hkvZrBMgFDi2Y/1AJee8auGK
8f7CAVsPqLiulZH1VszJoy/9+agjvBvbk+DpqROOjHCfA0JGQ9sGM4WEQ2iv5+z1ZS0QP+jM7beh
xyxaBFrKnwMeBZUBNOnkAODQiLwa3+VvMjP9hJgce1PTLhyjU3ytpYLPHasCmsdvcfeKK152EVek
z4mh6cAIdM0XzfMMFI3t72z6vTr8MsjsE4FGTA2l5sY2VySMFFavOMvnELWd8Pe3oDnuXPk6JAgf
2dRqX+sdaffKGjR9NQJuNP1NpV3jdk4WBrq9G2i3woKldRPJvHiTu8TJ3LBqfEXqjZJIx275T+k5
5axrBESUFTfm9mTxbrMVEj//mSHwPC82Qlv3jZEXJJ0pmw5QaPdXW1hsNvkGkctCouMBSKJD5tQh
0OlQEUcdzEAbMaQtt1RJ/+2VixuT+mkuO37EmSxWN0gCcScQHWtd58s6sG8OygGJ80iflhsMIjKc
2OwfyOhWSn77RFuQDs6II7ScSFfuphU122K1TCw3H93GRAHZj7fH+mSDdrC+h4l1dMbyDmBjTa06
8BfCfzChBXZBDjjTs/b96CYH+hlBNBxOfX3c8swVVMrLVuZvxKwFCdgVud49Xw49KoPS3qix68yg
U3zYvgm/wqEfp0OC95AYu+s4G8EBYEpl0KjG2J6gWqzvm2VwHnX9admdnA6AY6WA0WcOJY+k7+Ct
e8PVbnxv20H5MmaMfHtud18eLW0BldhuBSn5mYfqRqM0bYQAujrrIgPd93vwNhOa6bWgWtanxpX6
hpXPRBaEW5RlA5udye/OQbqzbdX9fnkYhvvhqr4Bpgr/QI8apYol8Ep4AuJa/pWQkpyUte4CcpFG
x15m3+ulhsBPKsj1sAuCBoH1hHMXzoKFx5R1wrypaznGTLMaHk9F8lgT/4+HyZL8eSz8T61+dhUt
0nQygHzSCX+PdwjaAkCZqF6HXjcYqnBRbyMDu9gRfxmErIF0kveZxZVXzLE+jrzhqAZjj+LDGvfW
PSFMv7/3DFt6JTs++qUTfXeisgYrfpWbfECpecMfonb+Xx+Mz5ICRn910XiQ27Xpq+bEJdXbwWnx
0JoAu6Zp4ouAiWRy0iFCsH9d9m3b6LUwjRbL+yq25ZgsQjLEncmI86NJ69SoYnUXK2Dw7GpaCPG4
jVwNDSThiUMGsPs5diM6x2lVXHyzxJRe/pBjlUuFbpFMn/lemwe/zgdiqj9OSHEQerwtsoX6ACs6
pcYMUZLxdhtZHjQ0bxZ6C8O+9lpjgMuvXr7HU7jnQQDvcMru6s67U3Uae1QTA6LLbWHyzDmclfMF
W44ygeN5ydXlB/KficFT2soWd2Gd8iPJb0w+jmcFmN4pzDeTAo1qPYo/UIVVIV2Q6eBcD8QDEeTe
Z8P9rYL0me/9MQLHTQNJV008QJ/fsDF8zp6kV7S63z26W7yqZwUE8NdqkzuMTHEUSYdOC9z1JwWL
qFUtsUrV+GmqGkhXtFlsVc3TyWp09RoVRQ57dhAKsi/EDLYmiG2esCHuxWHkpx8ktub0ZXNJ4GD2
aisr1VlvwcuIQqeCd7rNsxhYACoTmoEYtxcAiQ1uv9/XhyJkedkq1TBLZA8PuV82NOMOZJlULqxR
lfJIVc+0aWOLBzV7oih0MhL2odiBbfuDpgxeww7r9Oyf5fCAa/TZKQTckc2mtqfQHFfMxCcgdY5p
XawwOurroSAj2OxsirrTbDgRUEze2gNEAaxojzSVe2kuhkvdinSTxwMl/RWokBzZFeB8GTFHqnXo
ghdoh0tpM1Hl05jUYAnHhYGU//11H3WRh4tiA/vBf5V0BJvIHAv+KndzYSWCx8e0FQp6JXx6C6bk
TQVLMzmz85RLDJv5YwnLNsNaq6jZLsLukmupr3isAqB41cVS6F1E6SP8PtBlGP9jJzMZYiYslgP2
V0ob+WAz4gtJHGxSF8SYQZiXrVBaRW6z3i6j+uR3QucZHOgaPgbdKR10T83xAtb5D93B5muHfIAz
5ciM57urEbf3Z43V2g1QeCMkuQICU0HItVnjQzwxK+RZp5d4Wbz1smtisPATPdPE+8SCPvT/Mu1L
wQ7ma5fo5AQ5FYF2vOk5Wt/o/9C+MmxfQXVVVBUxrrZq7A4W2j2odC65skwdCyw0z1z38sMUsQ1j
uMlmEOyJRpLTxl3jkfhcYHHNr6OCZuyv2W+ZThIFDcOYfvm+HAVysXCku1Xuz8YAKQysrGRkUXx5
shn+xUo4EMYD3N6XFWcxYgCz/EON+VhfLJvVqs5/guY8FfO2Z8pQ4gUUvjyzFeoF90DrarCYiwFi
lGKlaMH/EJQPSOHaX0LuDxxbckZi/I8ro9tqUADDu9lVjAqnDOGdaHup3syq2SCHBciAfZiuBcAc
OfFikP9Yy9USCusS4ke3bZWzI41WmkUA5YnIkYyLqI0LUVgdHBFEVCESjjx0an4LlcV05k4/kc8/
t8njpQ+ULt6jiY61w2fiKXi4WBjgr6J1YnNLqn4K173StUNZhpRA/DWf9A4+uY80xB9HEVy9pf7H
AAtTm/xs3XTAp/4gRPOW/FTxTtnn9VrHSUczugZHrYry9EPzgPQWu3Lk/WrXry1qnhF8t6Ah27MC
gjM/1hC3D+652/mULrbJPHL2Br1u5K8BwqaAtXf0sJNv8ZLauq+Cou9o+HMwy2bwUH6+fzYwNowg
iHyBKnN8BIePmc57S8vYihjw+z8VVdORZ/SVtRxf/NqIEcGjgdq3YuoPrFUUyYi/UvdlCneh801K
J42h1A+nO49tCE3t6CTPCVAppVThYXmTsrkZGSEjeWEDw2KzFfpbVsR2MaWB32aQW12HL5O9t+Rz
Cn/eaIhzUOhIHeanqfYdFswT5sU5aM4woCKYTdy9NR34xGcyeVZ3t5AG+DgXB8JEXlIr0P863DUo
Uqh0omBSKV3RBIYBj2XmIJpF244TtivXZJADjr2l2bUfC6xQsGzeygb8kC9/x6+g1GGgBH5wBi9w
NxP0rzrXWq05Z9FqGcIw02L6YtsUlws9Tx+gqlzw9HXNCjeKSxh7X80q0VnyeowTg1L0T/jOiKoN
eToaOfp8/sjKerCFR9F4Zc8y5pM7EjhsR+6+65CYrDiKP4wUEeirmr6Be5TE2hhZP1yIOpUQkF7G
ajiLKXXhM3Jyken50OUHzORrtkRt8W3lvReURcvgxyYKvJPUm91I61lte5Pqkl+mcB6cY/LIzK+Z
4jDkfLJIfBW76FaIZXGRF4GvKAdsufEOWZQ8YgOEy2MhHcMQuj4G+S8pIXZORX/4Euf53XQ9ZCgC
/Yk/wgs69Aq2gcfTm5gRbmxhS2jFxiX67MG3MyjXK12EGKNtTSzPj3+Q2NxxE6QVXvxMmnu6u8XI
rAbDDDwwpE4Oh3EwulHPHXoMq4kyXMIW+dlfvXWnylJtFdh2RNgPwWdS1tOU560ixM21RS7R1tkU
N03ldJDR1N899lCUqzIwOflRLHSAY8Vh1onY4zHEzcmQYPXanZmjuT1PJPmlbB205euUTT/DMLoM
fTGhAeeLlgwm1G4r1ggwtRezIdkXHhvMSQFFrYPjZxtNajn+KNwu5aMJ+HDdRBCx5bjw/ImiuebI
VUZ7P2pfGxM66DLUoQCZ2ypcIgED4/1gokGM6pncB/g6/nA3hMROuBgT5hb3SwTDrA8iV9nlwn92
UmCqexPGNLIv3dJkytkd6sezvzVdoNUQIj0q9+iVg9QmPdaz5i+9nEUQXk3pvhdQcFA7blsksKqV
9wtbz+7+OwLYpDgyRggkOo27OFVJfKVgsBKsmWUfPy50Ik5/gYwD/rqQRrfiEV/nZTsVfSDzlk8q
Mqkek2+5ddDz0FoKTWWgXc18Ly7Oe7cNRRugTtQ0k0fjRJf4K5umM9HJDYWbuxXmXHbp58qGeBzX
5YAAYtiUM/aB1/eaPlB4dU9HgyxMSrVAd/sdQIyVsUaK2iL+FxX9shTwXEfRsBIYRGbRdOagbZoq
mPZ/vPpGTJSyyVug3yDpvA+7pLlbyF/8YZvHNxcs9Ksu1A3XOLPMh6j/UuYgC9APnilssPPIpHGW
9jjlZubrLboBAUgjhvIJq0roGqhq23cf+KNHDWi34EJB7Mb8xYXCF4RqCOdpO3zRpaLsP74YgEc8
+27PA5zK+w+gwvqoXvmzwjyp2tXJAoMs4gtiHmeXipwio9mKPw5n2i/PAxLLWNyO6lht0gGc7pY7
FJWxMlAd+5l7FrsQu+EECZF0lOCKJy+Kg+CQE7kxACinOiyo+/c2FIgwots7zJ8mEyRkeAmZ0Ohb
QMsdLPwi9wrT89sG1BZJZbS1qHKwfXDzEI+7QgJ67/REGX+VGKOOullNoG8E6PsQjbZdofdkO8It
i3Q1kxJQwHj6kduPXrM2V7aaHXjXCY0gzWICA0BaG9QOQV1xArqDMVVU168fdSBnHPyZeskDi8CN
DQ4Pi6wEnyq+6VWmRXrH3z4UeuN89gTyP9q/6QglLWJXiPkIH/aH2/JCDlTWfzMbEDw/UINnV/UH
PYCf1fT4jnYJxsFA24j9QjLaMn/GAXeyk0UgVEPJUiDcP2OLJCrKRgP8teWxtlO8nvQZ79DZEKkf
LlqT0yTD9lu2ZGLxqNOdEC4yUuJ2e2rd96HrVJsRjZo2oYB0aTN6ePnrmvs3Yn0OaC7DYEVMg8cu
FFSqWB/6N1P0llAkQdokUbQ3eV3Y4FKXIalHcYtTILC4DMCMRCewIBrMTeKAKdP5OQPdSxhFd8/1
+oCr60A3g6PaG441weSwktbMu4S7AtdgolVjfdBclMAC7bmp+2eQWXoqm92nxYVFjVVaBFf7qygK
Mm5ouIzVGZMMW8IMo7x0VfKzf6agYh3EznjqdJF3cdx+39UmQIfFyu792PY6E64wYixnLYnjcvV7
Lx5PV1awWQnJ+ACl/rXGgsc+xo4FbfYcVIManDt/Qd5vwjHhDaAZyTiu/sDgRo5DSUnNdWjLhd38
7iKBgCfnWrQWk4iMcgw1PCRl72oAB4dKun11InIWbk40DoNlegzD3D5LOS9HBljh/Vc0QqKs+evO
fgKkPufcC07NEG8NmiWXsKzhj31x0iLTegzs1/1xg58mqayq9RyGyrws7eCbF6GCBkoBtqYMGZgy
DfifRKPYprnyWm3YJuWQ4Dgvop5CAGUniotKSUBMm9nflpjqBP/PnDaCbr78t+7ye5cdtPauXXky
SExOOcnNLfV6vs2cWRoSZ06is8tjhDgtYtFINnU6OxG7kl8AbhyqRwJZaCxRNeY83OSAtbkBdjuE
AI+zQN76w3C0R0kNN0BIDAlPBuvyEtc3ROQ5IAj3ENn5coCX+kt0D1oKiZnJYsVqeDBJVyKxsC7Z
pkKNQqwfVz09/LfK7QN2o4FiXvcotVkNOq+r7Qg2srQH12aDfvCTWURMFXLdVGvRs00x2NWrMIhI
OSfieDw1CvfhdKhxLIiVi0GEv7mYavCVaFqawMz1vO+de9/j2jVixcC7mLKzbBsOXYR/VYDJlH5+
HNgwzMSZ4Fbh2RnbzoqKFcRYzew/0y4jy53FpgIcUfmoLmw86iF3VDmirCgNAzd7CvXdagXZ1UOC
JADyztZdqzLyW5o1UmYfakS6eBOu4RICvSWQ15q5r6B/4QdhfTYcm6aRxeTj6UvKEQTmHtFcjcsx
DTkTY+8TOvpUu28WUBKZqFAD69OxYJbx6WWtFtoG+sxqFCj6SMbPJ9tB4nw4kD8CN2H+DeAcICbB
clNWzxqxdaDHemHS0bEyy0DPjSCtFPqDg4dp/Vd4ob4k92SBLiUmLlg1+2ibNLq3lbGRZw275dB6
1PJdiIN15qjPJ29aEAh98AOQLCbn+f3l1XrPXrITEjBmjf+oevF2XmrWRUYbJIrCDNa7qlolrUGP
/pT6DVGacMMT6JleNVsTod2xUuQEC0rUaIxVpEH/87+Y3t6TFL5oklp4h+QsL+8A9K/nRsq14tp6
MuuZAq3+MxzoBPVAwLehdpBCF2sVoPivxHmscVighVmAkC5Aq5tHRAB0nW1KOqjpsY26PH+OYfuR
HjMm5uagbI/gC768+FyGjyfxJT9Fjh0oi2TaRGGYBjurJImDuUli9unDZ6ZJaneN6afguoQgBfE4
68NtQTUrl01mqc9y/qjk9LFBWd/jrHjI2MteO7g3h61gfoJVBwuCZab/4Gf0MrbzvTS4u8Vvm1YO
SQ4WgkPFArbOSIepDwFVreIaC647Z+WHNWSmMAxeYnPpzmr+234tiPvAjp1sa6EwROQDUScslHBU
z4J2gZU85bprzlm56KXcfzx5oEK41JuROPXcS7uy4B4KJFwCMAaLjSRQ+JBeqUHH78qoxU3C3ula
Yj5NhkcOmQqT2ukL2l0zauAobG2ACcwTiRSXg01OdDk4gdzOtLq1r1sWtjWdc3yHKEn8Oygd53Nl
5QOLF0tDvfEgxJyowgTnOzIdRJEvduJCoY/6M5vZTtVywD8g4PM/iesAnUlqYtMas5bNxSGJihuJ
pH9A81hmmJ0fcUyWWQWN/7oVbdt0w0z08u1841sy0dNnoarCosT4i8z5pWO5aI9ngd6FcHA3ih7O
XUxRkh8xtwYY8hYhQJW1FBSiYGIbpmg9IIpERFTjTPNHWkZK7+Vr3BpbRXZ46UywzQ8BUMqJi03A
fyRNI1gOjxFG15onWlsWczBAIP50jCFr6tpJWLf/S/aYTkojs6lHudQ/lYliiI/XCeIsSuj5JOXr
mhAVOUG+z0wXkSLfaiBWaobAzIFHWadczYm0zNRw6Ez0VreqkCMAh338a0NtkZ+7IzdNQVpcnSda
MP8Gl0ivOiKu+A1i6KR2L7dQVBjKD2qgaGdm4UvaPVOLhcPrODF3zK2G0kRhHEy7iSO6k5wpsNih
f1ksEjOE5FlOjXNPNzOYdw0Nd2tqCI2H6cbnDf1Vk0tarTCJ+IhxTgMba0Hx/xTXON2gLyHkGzE5
0OIM3E2XtGnaObh+abEavS8+NU39OHepxvVq8pGkGcujJ4CtdgYJPQaXKl6bhN1Wy2j9+eWTCqd0
BuFLboQhCHM7lkDUf1shkmxxXvXOxFMdSmDtQznKAvulh4lq32GeVdPAX7SaoC2+L7b5g45LnQ/H
+vE7vULALa/t/ekjgyurDKv99tAZ8nRGBcCbkbZwVUjS9AnKSL16yDjEJctREVfwALSwglEypAYo
RYF5x0Pp5ctRn/RKS3AT6/SC0+U2AmwZOK5IVE697awQyjMVaa2VjmAG3X1GM292rO0MHeu+YG3m
cuy9QUKUE5Vftku7s77d9XEN+P+gfCtlo9zrkNGGR5qdKF+j5z0mfrzpo5cpFB0qFH8nZuFpyxXD
Tz1W3RJnDQbk+lol1TEAov1NeSjA23PEJL9FMhMKXBsgBj54Cbf7q/jOwLquA8NuggOJsMv0b7tC
KSWV1nqLT+vLrW6ShxBd1DlVv2QJ3LPYctIGaDr64u78ItqTKDqjRsgH3lHEAts1oYk5lEAE+bE4
I8LftNaQ8yDRZ2hAMHrYXr8vbyih/358+9ft/wlPfQQWcY/YaeeVkwezEjOwX8J23DMc05OGYGls
Hac8acPB444nJMfYpclDCr11C6NFeqYMuvsJLLC54NQ1Q4nbc0+zJrYFfpcWw+ZpGCqQPo28Byka
RYZnw3ilfU4ETV1CwTLTSlqhQl1Zufc/UJe7ux+fRB4ZDZrCHdkwZbvtacrpPGLeKzPR/6WaXHuC
8uyT2VP70ZWBPnr7tttCYlln2ZdWOa+BYY2/E+y1spJS9LLdISCFaWwHIyMs29UuKOJGX9IisfaG
bu2gnDVmgcc6BT8WAeyMAsl/bQOqrG30YpeYEmNIk3sG/yGU3+kWzmyy8SBIReKyqEj4ROeR24af
+NvEVhfyu8W84oytMMd+4qUgzX/0Bh6j1M3WKcS4HF85TGovg5PhFvn3tITTbvwOuJdSLtTQmgcQ
9rI3/1OAYt4kdC4oborebK6cBMb8Save1QDlD1HmxPs07QnJEo8lWm/9Voo4G4HJiaCZZIQrlgqk
1+pcHvlh6JJV+m3QrLsyn3UtmBWhggXUcjMblMZlHz7kAV9Xh3t5lNaBe+gQ7SuVAXHHvvAAcS9k
mx8TXCG91udbiT8dmDdjjVD4vwqNs99He81npOsazX+zAyGd8jVXa1DVesnzJtxiQ7z61ajQ9XkW
fOPXEXG4jMQ/gqGYKy4+93y80khJD1Nli2QOYGZVYmzDKIk3oAIO72MbNUptS81ccSCmVBwsfJWW
hde9JWiczMBa+QLSzarvNPzIpKEjUbmaG3DOM+DRAl2d/aBlmQPDkJEFs5rJ14pZ1Wfx0ubzL237
SQaEnU8rKu2gE951QiXZ1CHTCCqhgdMvovIxj9f50k+NIN/1XDpsyg9tI7+l8p7syOxc4yr5d5qa
b/XMSGRdHy3aeqXPp7PiCpp7yxi4ThO4dTOV+0xRwyrAjbab5P3dFNKh2tZrceHXkqldzg5oNXpN
Ybo7AZTwn1QQFAtpU3OQIgyG4gxTGtWCgir29MR4PIcT5DizzMrDy7L7Vc5d6+Rf96KS4/pCWFX8
wi8CJNtO+M3QCepeAyzUz+Rs2qTYbXYv+v/YAqhYeT8SaCyf6ciqvM09wRULPi7UNrTj4X4xlkUL
9RIua0+Ibd8TAVuUwfLl6mF0wGSoycS0EK/xk7XfvMo1piGJMAuUosxFECx1kiSwwktHfS2viLuR
EOf8Ym7ay4ENojx37O57wHsZ5xjqiruOS/gczycnYlNPkJzaidC/EDpNUhHdajksRf1mZXYP07o8
wYA4sfe6kMl9/agmq+AAQ25+QcNTbellHOIIMd3u+murQKfJXq/v9BdK2z5NzAxPNG++ztMkAS/H
qONDZqJ8te9GiDEfVkHGP0icU3AXH2fCfKgHLflE6JDEBkYBMn/HpRQVoNzlR7Jlu9NtDBEoMI5u
GJKjHhLaWIv8rTtMU+TWiFWtMDQFSUlyDmAo0W505B9+MpuRZhYT3BHiQvBABFRP9Szmd2LYH4wV
L1r0WT5l6y6FlyDNCkidMnVPhoHTO7ghhXbYeY/h9hrT3kVZ+TE1jnQ9lxX5qn8CGSb6kCLojiKP
583V7+nt2flqsf/Tdj+fk5UR7zWYy9+oaN2xT0fyr6sTkpi/CX/2ukiRM7Mkd2ShjGZ3vvELuV2v
7j5psvR4vs665nrnUXymMs5Ox1d3fU73t2pJOaux3EidEcksU/heTRjd9FHZ3BfR/Or08l2i1TNa
eFuz0ejDxYO1jACGHD+grGBGGeUDi5f676B8wBnjEoN1LuXgG7FDFhrGCnhaeKqMXcSByJ0pobMt
y86NDq7rpO9EdwinyelSUjakuFzdVjkfR7fmvbbV1OtbLUKdPS9kg74ZQyh4i0IJigAwH40bmu9a
Clj7BUJCdc4ByUE2GFekPBgcSBMK3vsNqK4CbkIAYtHYKcW6pF268vqSVMcqbRA/Mxd5iKPkTewI
8cBdUNPOib+w2AbkfS+cPM+f9qUPANiI9U5H0VQjqkhstuN5NmrDtvkP2pI/rVWwUqZGfs1OXKSx
KW5hpjnUm7VC/uXgagP6vBiEjpj7cf3bb45PIvu/LEH+bH/oPcEqXH9cBNZ3IoGlSRs4s55PTUDN
w6KB4mC4la0sNNw42W2HW+Y5xIfYwTdvIvCqx5kvPcogzmr3Cnv4et19Qo+/sZEjUBFxHe0STd0N
Hryj1bZJTeXb4iRtUn7f52f19d9gaswo3+P4dBM2Lxbx6aZt5yhJMXUSXRwWztC/vQM5xeaMiylV
7LdZyULEp15Zm9Ey/OOT5UjgMH2QwAwA8wfcJB7GXx2ro3tZO6otimcCQ1nuaOv8+458zY4VQwrt
lIu9/ERO+mlgzTwXSK+HItvc/hyK6lCVs7226CTmytm1sGi7GHARkqMAZqpBgEzK2EYLiQ6mBDoU
icfd6M7IHEbEpc4WBlYElseLiQr7jxtSuyj8xRyDssgqmyu0r7KMWZHJbfVJBDqhLnyRjpsUHR8R
m/w9Ngci5DVEozr73n3Y4d0fgQL+Cxfx2V4mOeAmqhBcFB9rfkyKkDtYzqc6N7MVpLVzjQhIziZr
2DqnmGFnwa6gUc0ID/isKBNPOIg0N5VB148hV9gC3o6qNn5Ecb2twnaQg8nhzswqAmXXP3/MZD+2
BTyUFHGRjvGRiDfPwukCBRhrnPgSM1H6VKBqAEDVqjVrJBBEtQZqMf34EWUEQ7hWYIpsp9PTjt0W
OmBvVl9pDiv0j5arprxBRHi96oU1iXFu+GrSR1bs7yj8nE0TGxu7VktT8cgL+Vg6SNoLU/8wvnKM
Bu1aVgSM1f/q26+36zi+gQxkKHiVc8Dpan6hsIff3vf7fRLOX0XGm4eWfIUMDUseo+rWQcJxhbg+
y3oLMJWA27TmGWnUZRLYuwCg/nLEfK7gqoWlopczgHM+Swk6e/1sroM8jQj3EYcZLr4eoJY469f+
hczdGLGKhvPEc/EuA0j4k6vnHgHyJWeK5eIElvkBkDA7bpZfOKF2ROoRG6+XsDB8ekz8mFyzWe6o
EM6qEhHu2gz/qy2mq1ej/8KxuIn7vmRuOJkGJ5aGrdWTKtkQG1Z7wLbLgmgV7JhLhU0trY5hKe7B
VZFSaMGEVRnUrDwxLZ8Yv4SBfIkTzh+RaTcOjWZVs/vQKXDsnyzevTScw39cx0jdA8REn806RBMi
kWyESGKEC2SyR7QuYQZ/9uYwkUsJqPdtCXgsi2AO5vEEXWvRJ/Sshjc05DvrPxtFq7O99rsFNpRs
jrSnsKufg6cNGGb6vfWoQ7gXe/EFWBQoCkuNFQPzs5F8mSzypXF/NhcKOoYPsPonUw0vliWY3/M0
gY8MU7gU0lesyZTQPoV6arQBqY49f0ydD1O/OxonW+MdgAjpn4iRQw6sApvOBQDtTCSZTxPfPRwV
Y8eRY+0xTbwS4OkUKzWyO7+H6VeeK7OJWVK1SncJRmkzBTNRkG6MYcMa5+tLRikuh/Rg94sSOp4o
QeSpaX0Z3hxdSiSqyQiU7jjJFOukQLwCGsBj7r2my9d6x9E8RHjF0tlpE9NoHRxrY7RZ/OSlIP9J
yh64YXznaOB3HgI2plyJTz9gsszmA+iOHHqpc4Lg0f3+ipmjpzoAu0w+50UX3JjD+OPXiax2E5+T
+Dy9W9UDPQ/YiDp3rK1x9cKBSa73jNkKSfU+iCsRqoh+aNgzz4nks8pGgsPFnN5AU2NWttDosWVT
bywbSGppZQH106wbDU5ZM/CZBTfzFnMbwsozkdBXqEBHgo8O2AqZHa3GvE7tG/ooyv2pz21lbUkE
J+InO35y9a3WTYc5zBv+1/B0W08GTc30UmtVvPebWl237fjO7nkxsb3uGFiY9aOP/t4FBxvoujl/
eqdJpwjiIigBuVuKJKHoOKLgLaX2I6jW82BTmekqt+vWXzmodciBWU/azhO5fuRFlHX1ehBqTiEB
9mGWnOUTHFQekzM3UQSaw5hI7e8/RMIKS/Sdn5oVkt38pZQS+/b8N6Iahy4GzTlalpc+PK87qyph
3s+nPN5iudkNDwQ1t/Ewv8KI3pqXAJGfwlgq2uriTaRRl5/dczViQU+KWLGgEL2ZGrbdxG6ibkzY
oxoIlEd010PQ1KvJjZIJoFTB294G5D63KQkituWGbKz8G3w48SBa9QetkUpwoyLczH4NrwnqCTmC
VYuZG6cG6loAfX/D7m+gO/EqDKbissqLFvR7HdJQ5sE9iB2/IkAeu0gW0IhoZB03BujAYqugB/VH
E41pLs/JJQR8ya50RRgMOWJFK5g+WQ2ecwu7ydDtNpMf1HSw3plrmxKjk0FJlKMoC7aEYqE6n6rK
Fse/xUopyTpLlG1LrZMfNjgMW3zq1UBJ/BlyEytCk3VqbLC9MhBtxIc725xGWoG4tRihrZvPmNlL
3fwLVbX8jUB8Tzhvfnwrc6P8j3IEnqJCghyBCL9b8u8qtt4ld+FRHgxgf9WPpY8Uti/MfSP++RdX
Y3bRJFROsdZPaZA+u8F1gajX5oskkfaHIBsCVMlbnWNGn3F7woTf/jHpKRvgILVblQPaHE9GW3Oj
8oY2ipW4jeMNh8B36+UBeNCQ4d92hzLhE5p97TTYor93yW3J0EH02DjkNfu1EfjXxmKt5/PD0bZF
CYPJgufP3AwExBGnS+Qz52cadF1kTIIM/n+qqeH9XoRMCt0+YGcs3zbmq1fM/mfHgF05z6feIs3z
NUkFuElVG+lG906maQ5VDx+nXc/WcyJbW29RVGEQTMgA4s8cs7Rt4Z/BHHR/pnOEqOgUhrOv5jMM
ISUES7986yXEAd6UUKiREMCQaLJ+dsC1P4xoFyy6fJgtNze2oxMZAlp75r0kOlgIe2ZbmpGykZYu
axGX/Z7YVgGJ25YbFy7aHpwlZs1SXNsivfvTLE0k14VnItBj8bmnvZitKi+1wuDGcVkFuU0CtDXU
Gj+YWMK/pXa1tv6hXcDChHCiMVBWNzGSeZBMdaLkBOHtCOkdyXhCTc8sagRP44grDz42Jd+1z/t0
x6GxQRDKBgYC6iO+mHC4bxqwVDWkgE2xm1FbP1yPj1WNxqZIJGdP98JvBEch8zw732rj9txsvWzj
W0GqyYNS25gYkbJekXFK5rbKYjpn4OWhZChmIJRhSI5KFT1x2NQSPE6wVo6ixnyM64ZkhEAL/fwC
YczD8USnsjPmrLuUTSVR2DkFGxU6Zax7bkAJ9r7nW3nnFXDKIxeLHHaZ9Mkt4CASr2qGJNUCwvp5
AvPpTYJYSfsmBi7WeluDjIColcsVyGFNck9ubnxJuaVPB/pnLQ3qHHIcVuSHn4ICyYhAYz6Dp0ma
Q5NXeawbURQ96uY4akRzNHIB07UMnsujAOqAKekyPQSYVMoSrHimetT/hGTEDb8oW4/M8647nD5h
y7Trsc8KD6geg3iQu+U5m4fPfKwbhrz0FZxIcR+cksbTDU8sV6uSSyIs39NC04xDeHACdzSgT1ba
qOKkuCZT9lkNJdkCznd7wWN3RkFab+n8/UxmnAK8MlyY0bGZurbG7hCNMyVwfsRHUviLVQQOitK5
HVDilORjpJVFgSjS6hV/xLtrMgYj+a6YYOzU3B0S7TRSj5yjtjMFKNqp9izIA3SjhXLzrql0oSpD
NKXZCOzMkeHQz5UQIoAC0HIcF8IQtyx7f1eBwYHcepPgjF7rRL2+2FYXp3BBmbspq30Bq4Mgay0O
HuylOmtjBPJd0Gm9l8ab/zR+eYFRKkRXM5JLniLsKv9Pl15kTTXrPuLwUkpQvs6rdJUZ+g6CEjlb
GB7iG4qXRXhUmWSrF6HQ5r1I47+QUeVHBy1jUrlB92JFGTY/Vg6vY1WoKIpB8szaBykUie4ZapB9
15gy8heECxyvBlJhrGifwOHvDxXypwhQfO4lu5Hqe/V3sHqvSV6mHTStE1oGq0taZnzhZ+sMg6Rl
owl1Yr6S80GB+gjIpChLd8L5Ky8YTdMohYc4oVBALAzVdVy3jP533qutH4liWU0Yg2V+ldtnEb90
D53vkN0voKPxcnsSlNt4hZX2WwGf/Vpce5y3EcxMG7Ef6HijYKy4dNFh5dZsJjv4PzOfU8wb1vUy
F/as1KNrZxVuIlMJEipCVYoZUlbO8pu7u6DlAcCa3DgkA4HVnQlRaQ4Z+W2V9KGAXxIPedzPMGGQ
Tu4ZHDQWuxu8W0LNcYr8uN/bIpvquPJfFDRhg2W5zNTG+xRmS7O+HkwNFpgYuhr9U3/Ra5YFL3BD
8sSw6sIu8ywoyWVVSpFKjEPjy4L7LdYOWbihQUcQV+Rpah98/gNrxvnaW7/THwTQdaJPZpK8Z+Sl
0qbYxjxQYzoDxSJaPOOdkYCtM6MnJk2uoPK5x42PmQ+KFfDYZ7hjhlOLbVZlwoLQASSd7bJPaKgF
geqhsXNHtJrlblKDKaYhLFS+aNwSJdYnFyBHr6qRgdmLXlHbqq5+XOBfV2svV/YFQJm2LfJ9H0M7
6BDnZEDDN7PEu7gzRypgcq52AQ1fkM8n6TZEPFiogBblitUVTsP4k8C8MSSW6vb6zflwriJx23mx
Qq1oWB8Dy+aLztSsmuM+M16MR3ck/zJPNGxBClqCwBVE4P3M5+B9/LP6wunxk1egurFnNck8AwNq
wKfds+RKoZEhS3bx6BMGjlvwq8DeFzdDKtMGMoKfhgBRSqvqI/3+yXDtRIKiFWbVCLqi97S7sE74
gXUWBJ446uMBeE/N4fVktYcaFyvcHXEmsuBLpdMPCC30xeKEEE4nWpJxKEihEXdIwHwDRXr22Ggi
+bB02JQTTRQkTmka0Ci3IUXBbYRFifNwiHJPVTznik4jz+rCQ+IgLkwM0+0ZbeigLbi98vLPxKPI
UGCHNhjplVR8IKjcXsAmdITom6tJ2tG5FZKOtc+CP1/EHdTskpY73abnbXlaLTOpGBvgK1GGgl/K
gOUI7Ke0nkH6Xtl7pqyByOsnAOBvn/UMSJIeiPhH4anxj3SJOcVe/IcETcgC5EIVuh7p9gnz85Z/
5w+1n50yyxdusDyp20CXLMQuLxqBr5ljBnKzUeusaNLSksHzt/zqCZxX3Ddwkx1HU771ZF7k3hXL
2O+IHVEaIsqzF2IvggoH6jOANfxFhv/M8v+F/uYrn1eCzOUHa0NwXOLXPswrAFMfZVomtQK3rVQR
101HZH0z0+cvMK40oU2BWfJo3vzfTnMz7dzZhO06amZ/ASU7yV73zhUvdwM8JOz1lbHjkW/ZLFEi
+9LWLT9ykp33SnPHABETnqQn1E4F6VtJ3glOZLFD4l6Zzj1euJbstf9fdJRbGn99+Rzk/Cs36P97
qMkmPjuHEwyLnN/lJnEM+9M0k91qbHeeCpusiPxvpUnzq2dhZp5kUwah7435LOFkJ14bAYoc6C7M
ZePEPupgNjF2OkePsdvE1f2ZAfiYgs9QKg04lI28IUMAEPKkkSr1cE5sYEbd/4XRp3FDYBArxZfC
mmmls3Xru7HvvBtoBUPgwb6IhxDWEI4eaIoukYvojSadkQgtsR9m01RqJck3YNd5Q6nKgoxVCvDC
WdQSNRpxWKoAA0+ImVtLxYBDLI4a6u2fYJYoLlf5ge5IR81pHahabMh3OJ7OSRTAznLSSES13cJp
uycgSUpgmR1wVlcNtAKy6NIc34eSqdTFGH4i1arJmDcaXo6pHFDJ0guUQhaIRHUfQJjr3HCa/xNe
zu6WF3z/TQc/GLreIJ5/reLFGzHUuYhSyD/AU24ovsOgTuw8f1dx1S27JY1b6UxJkbZlsYrQU+PC
jfJeKic1mQT7bdMdIw7Ch1oyrdTjOZQAIC15PozyltV7kTSsSK+6BbwSDmdckdaZZUgIV+H5c9L1
r8TIrGef9JsA5slH3rSXSyDpyW6PS/kwKesx3ohHL3YFtQTw7tu61k32bA48NYRrShOFUhK54EEr
UGjSNji/YkTMS+VrxiQpgnI+XCfl515yGOM9Q5qWUIic4GBdWJvN2XxttKIx5ivk9s2xIMC2UBUM
BnqsYV8+7pp4Jjxm2BmrdkbtIo3BSExDMZedT7T+GXEM3IO9xMRh/wGH6ohJltyx8/U+V5ws1M4B
xV+yzwV9+5BBCDDnQi8ztvk0sp4k/e4eBUGoXKWWe8Y02Hr43KgnzZDCED63AC0UstrtEp/5MsXt
U6LhKBoZDiK/TqWCNvT2AXIe7s8qbkfqZfR5cd0gpN3ZD8xrw+CatAIrt8hw4bEsQOQyF5obJhpU
vZWGZPukFCJ2dZRAooe7RCry1tI5Wyet9/a/cuXl4ipdFd2BtoWYIbxoAXGnTfF+WH+CJNBa3HMF
KCbRM/3Ak5e7KeC3A9CmEhaFxsvSJFbyjx5ln67EDHI6ICfyD7U40TFO3w91tuRn/OIxH9ofZwrD
LGhIl0WROLnvsgQZve7ENIjWbnfImr1L8ZNAx9pHjmwT7LUOihxx1G/xzLnk5E6ERKrl0W0nDP/q
1dIWPDeZrZrt4S+dIHnvPDubbkhiEi0Z7AqswjkVe+vFJ6tFqoYU1iUFQDj8pEtpKB9l+S6vSL4Q
ccd874OqyhmnKRkD8xDWBg6ZIXkrDEsIR0jnOledevLQBaUYkqduiz4I12sXfNvw4ZT39AoaJa7o
jc2rUWr6I/gdBrRNgmgPCSDG86ELTh/mGd1yY2tuBKRVhB0nhqEe07ivDYIQkOONPc1ZX/lCAZRr
E7ea9SdCnajxYpq3zYRzBxhox8TuwJJ7L8mB0iqzjxIRjAc4IQxORuyMkElSobvD+9GPC8vlZA9F
ePMkawwIrrEyoy2Kwq4VbcNzGVTHupwyJmandsJCudzm0PylsDTkq8A6RweFc0l0xc0jaSSbnY+S
w8mK+UGHd9Hfq9Nti3kK25EcclP1IMxDPfvVi2PFnd7aclKPN6gD2eYxA7gewhtwPrxVi3+pOgJ6
cr0VDdLcRJMvUzAhbwmD2wG5yi3iJrPQPxPIJu6DeN+WISDAOKe1u/RGrs35BjOM1FVsfOWNdCnI
IHogOzhZLBd5KL/TkmVoCNFs84mI7CnkvFLfZ/CMF5RFZcWNj2r5sce94DM/u2Htcd1VVg2tglRb
wjCKBnkTVaNvoxQjwGYSyin5u20u1MGmHtMlE4koNsHQ32U3TTYUwpxxGnYD2BBNfWabRouha86/
XNy5ieGZw2WK/E6DqgwJJ+VznYeYDJQSjAi0o1EH+cWp9FI+6BQXZIfTwDRPLD6DV4nyUFPZcpoa
MDL83ZhHZn77OsRBsLel2MhI+4l1XRSp4tbR2fsZ7y1148BvRLtcV9GcoPESufSbGBYnUSZbHxIZ
BwVpRYm2fKPjZzsQCjiXTbYU3FYMdXQB3RfdX9M7rcDEZ3T7fm6mGlnDnZKUAQnGiaF76+qP6iJo
/JMbJEMcqj/aF1l9G9sglh6WT8YfHtn3+ITzXCrjNhWsE3074XGzROIZ0haTh8T2ARbGSXpkp4d8
JGPAVa3amg6+SOWAluV3J8i40a/dXOvNIV8ur2CR8nBPwM+G0bqGt1xiLIlhC821BzfytcKiCTEr
kyazX1A1AW4+KqonLFAnjfkhb50yYCUwPJJcE1zue3KL50F/S0NyKLwi8EQC56cyKv/OdVXZ1iBN
C9A14iP/L3NrLLIaUIQpyumxrmQZI5Fb1SNSvOkd730O8tkQWVzlo+y+w2SoKkoLvCo0k6GtZnE6
W+R3/YENlVHwgKWgm7SzGRRTBVDtihUhkUL+QCjSsFJEwSacOO3Kir6WqLiBwzhNs0RGALqbO9Il
cx/oS91yzNbpg5CLhvVGUig3RX67ZOE82/OcY3sI5YOGLq/FHjWjtXeqAYsbT8tbf07d2Jkv3UY/
lDVk/E303bcu2KzrkbaALJqozfgsnnZ4yXC2NdDnoITmEX9cH56gfBg5mnvBSllq/vMd7zQfF9q2
9mlQi7/HMefYRibjLa8kAH69KDcmBpy7AyEvyLR+T7KNhC31sIVx9crXWSs3kE/UjVknb9/orq3P
CQLAkuPf0KkVjjykoiqjZZjOS8DGlwVp33FRL6MPNFJexn6BYZ6f7c0IlVAnjh+IbFa4FT8BHW5z
2OqX5J2KME/nswHUfN1tH824e55OJj3/iBKLDyQA1ix8+tq8l6P8gDn2vsNNScXrBW+nBudgZOAm
fHpijqR8s/8eceUh20JjjtqoaoKYi+PsAMVTWQ3w1mW5IY35IFookOvTiN7FPuslQa7VtVns/KUe
5TnH/SF71XKWAWhFNhQTDbo2vC6qSE4951d0W4ejwB78vugcl4lCPT4d0Bn6nDAd+IPaebcKYApr
tCz7iVhZVN4/Eh0wwrBC2+R8ZgO5rXJM3Ah+JvBpYgUoeBtj4eOiHZzzerxen9shBgmmoc0VsCxg
1BCGncgR10ex8GyBsBA5wu1N8pJimhANUHtAYgnzVJt5bxI6cDkNCYZRgY4wdXfGrLgtg4CIzHod
Dau04tTNsWn7wZwpJ7HYq4l7MqA3rJGIBVymupCTM+XkX6qgE5vTJh60bblLQdfmSbhSHLWD1yRn
rEaL3YGS0B+mieZ4AWdFFBiYWxrjRF0B363xlakypgdO1v/OmaKtYLV/jO6x3mr6KiH9hCo/18L3
BsgooTnKFlzpKoK/n3XEAalfZJwSbwVlXRWLeY1AGxNHmrc1awV/h2sxY7K/uAZXSISBsCatAEn9
VJyMI6fiuFLUH0ITaCeI6fHqis4g+3ZXoA/ShH6XeF4aBrJoivcGNmsAzK/u2Mo8mAiPiTxBNn6i
zWCORSkiuTqUZtb3tqcSUJ3DTwP9WezqniyP2vCKQHA8321lwu0hvpCPzIx3fUP1z1R9laCp0Csw
vRffS8Bi9AiszQpvVSClJS4XWGJhoQYYQ0YzzlcjbEYwlPsrCV4gVU5vZPL3s0nLP769UHd0auE6
xdsuJEHsQXebJ1R9vTAbQfZGHTQXb0WUrAGyTqJTYcppLUPilCITL8TFoQQwNhLkxlO2IdtdD8Us
q3VZP3OvwacmIkwvgdDcpYBVAjPoOVgStLymB8Ifn47Tw4a0ZdWCRs8dHZXANHb4ns8N6tOKhOU7
ztwjTuz2VO9or8DFGE+LIhb4dVxBKuaWGleVjgrA9Aj8zysgF9dhTjPgjRPvqPd1iD8L4RqilxbC
0+cKXQggsg5dTn6r8BMcZLKYyy4uY/H2ZW0kRSSAqsylmn9mj3jSjyGSlj+E/ST3V4vMUppVE6CB
KhZq/S1qX1nno38Ux76y+cRt1uwXTe3Kuke/cA/p1H2lEZZz9wrt2PNzcVwOprzEgGxxwKcq5gpl
sdqLkrTt+lQohjWVNPRo7Xy/Q13Mlg+KNtH/kelTvY1n8COwuMzmkZ5oJKgJL+eu7wnbVPbOQ0Ch
i4MFuyP1bg2FEiXrLoDcdrUoY04IbG3hW/P4+VqJTzMmfee0hZf9a+Nl6fzqa/llkFZPBN3syFtC
n51jOWz0zLU5UpZJT+/fJOitu4N9dSAUgd97+Sl7N2VxTNARWTzCSi7FSq730S4o+B3Y5E3I+i+8
XRfLu55EzewtSTO1XoTdtZpv0hLqfgE8kMnHHB/xm3h+H712rrbnhhY4gbEoCVN7wXSbjjMrVnmJ
5xt1kUxz6NyzMRNV+DAfsTzR/Q2pxzu2AR/tN2eIP2UJUZIGgj3kKudAKUfom2B/vZPdVK5Vuoub
4s33P3A3CcvzvHN7Skd9N1v280IGVD7HT6mKJSGEdoYNkdhiueCO/OMbWyIc04IF0FCgu3J5RYm1
f9FyI43nGXezKio0/oSvi9dHjEfAuTG49mh1MUhjdOsY7fs6z9pbAzCrVbB72HSF+Kq4NZ5en80b
+Tj2myKyYsm87fE6YIY8HdtAM3ig6P0GxbdwiVTa33RbPNE1aU2zZU5ywQf/qiT4+K30N/Yma3TH
WCC+JNH5CJLnNQZL9MuV9fMs5mCUqYfkl/EZ9g2vDRKYoOR7wu/UFMx153XIxSt8gxLoEXzRuH//
BblWP24zNEHJe6mwyyCXXU55rQLkoOXM78D79audnfgNRGVYh+z3KCA4VyuIRv/x+lwN7JKG9hut
qhmwQeWmTFYD7EHN+R6gJpC3l44VeqoytwFVb1kSfddN6zqtLgGXdTcRyfJtbrG3z4DNv4CSpbO/
alS1o3Jacg3pWnH5vtP/NU8eWkCl9JEtsit0uCmU51XsKSsy/umgauKKUjQBizkGID7SAudd0DTw
rlvM6GxOfZkBqBoVtcRnqnvq1ddGvM2dnqe9vOrr2+QFPhjhlOAVN6vnC2Xb8VK56pr4PlyrIhDZ
iYEuesI5MLGn+Z3/Jzq8z6xtZiNVE+K9yrFoGZ9UIMkdct4VA2Avq2MWv6gJfLzrAiXbkeGIVSoA
eZoK4BgMs5Ui1+NoW5Y/EdP87hGdy5mY8RHJvSdcmX9Fobt8UO5/hAF+WGdPdLBRUIITbicZSkkM
38PVPaTXuF0q/cJmGtDLNb8a2bCgyugGLqrAdiANRUv4d2DQQKgOuCj0Dzh2tJm7NGyeqUGJ3TkB
2QN1jxY11YOSzhrVKx7/wQ4iuYkOloBTujtoToxCIe4tYg8i5UpFLgiLqZ2PxojpQBzuYXCs7YW5
0oLfEUQafDAywGWqO40WPufa1Ix0ysXYBthH+gLkbO5fB7PAmrlp4GLF4eOwwN6D2f4ySRpEwno0
5w6bUbgn3dC69Mdq93auFCwhETdANQOSbN34vYUmlKtwx3uivkBK7747DDtsOocuQaRx2Mt2VVan
7Tt8kwFTtFNLgdEtUzTC+56M7tiBhLuMKwr/dsL7cXPUkk3N1GXJcfYOugcB9Hfcc6uAQ9zk5LPT
omNSZAKZUQ1KF5P2mQ3xAIzgNQTzIMOndxqJUMKBjUFPtU773l4Y1ntGpodnq3/exSGRxX8ktfcU
B2sWEItHHkvaYYWTWRtVg3ihKX3kJCDPpb02s3Zo3e/eiwU4rzgU4a3KU6/nrcYPEnfo7QF2mohx
ACPfbIUd/wQSkrWG5J6Id5qYy1K3h460eKRqO6IRLWOR02/nk9x4Z4+Y4prd7EDiSoUJQInWjT6H
6G2OzrxE48WA3WKbUoUm23q+l0bFnf28mJ2BaTjTL7o6UMiTlRsZ9uerwh4miJ5w8EBAsGMfs8a8
wLhE7PsodMGoyivIcqdlpNNO/uM2TN0rm+jn1UjyJzSsaYN/X/gcx/YDasZGdEK8cpz1pURZHp3d
F+95/DM0j68ijrEdh2ULxxOwiwgKiIx15xdVVwaq7vLQUz4QsLHipwXgU4ASfoAAMvBapPoegKRA
Q3WBE5rrzoycNlZJlbndoua+Y0Q91XDle6g7W7onWtixaJU4j1cJcIWZDGmBTNaZX4QquPx+kLRb
AJGdr9kdS/6MzYVAA3PfIp0mird1Lhiu7SzbR4xNnj9XBjfsl+tmJ1JKBlXKbtsD6tAe2/joO8pi
534zPalTkcj+32BAi6jKMmnPdz1VZkxHPMfvHIJ74pvBwZBNTJhaO8IT4jxDejNoySZTwkrBBBvh
Q93x7t+syvyRcCia/3vH9VngORvh2qmALoIz0ZTegopNHfsQMA9xUk4tnTLP7T5FCnpKiq/yqSmT
Dc+XRyIWVkims49gjwp5ZD2RfQbJSr0rQm5e8z0K+UFAuF5xNA/lsPqPZVE+hZzToZpJA85DJrPP
PRLM+IfZNLpzXw0hsYn0WIfPu2ckkqFsDba5yPS+fRq4TMrfM99dRqxvief32OHqpyr6YIVj88/S
AFtk7/bFNDKpYpJAcBWaRm89awOhO4DyfL9fRr2QToNOaKEWbDM2qwqNnGG1rYkkk+ePuCi4InI8
9LZFqUviwesPVT6RQgcjMTzVN2MYbjqj93rPJili/vdzd5rCSXt/VkR398WLSkisMXemL39XbOfT
yO9L2tShqRK/6EQS6vqT9VF5zceVV6DdIur0v/Fo/deGxMRTAuWNhL1XdguF20czbFcUk3moc/7y
GApUhAj6jQKRaqY/6gvOCOQRC3RRZ5FTz1QPE1DOUWp8zwbNgECh2ONf34xe041soNy6we8m6ld9
+sK+6+W9bbLEM6ltLYKcnfa9bG3LgFNa3UD7+3zVRuN0mR2S/5FWe6dqpS8JEKafUOUckls9PyQq
ef7a3bfora/W3UZtul2cJX/NBoDCV9HNgfmqdMHdwhwRfZnoAx5WewJtIyjWZ2rB1zwrRKFmrTQR
dcZh0R5fYQCb9D7xYZMzzPH4wpa0w5fWApzI4EtDU80FJX3Y4osJTODXmxAfvOnxpfv0f0uwmWJR
/A2cWQI1ecktYujPXEoO58VnSayeD3fgKvDyJbCK2TZjDrlMwE+kV0l6jkIQvlEXvaAbfDj84vtN
6n4HN8t+VAyvRLYrwW8Mgv0Vd2bv2wcGTox6+tGmPmz0daDDEBIPgz050muyE7WF5Qw90aB2cc2q
HUbWa9BPk+mLMPXUgb54c5AIRWN7a649umGcJy85eSmpi6fdXpihwSIcFQdZdmeG9Anp6lrxgqkg
7Z843tsWOzeppN/AymNGjqhrvCPf+l255nuJcm3ZijatJTgT9Yh4FdlpSVvP3RNoegAuxaF1UFhK
ca+rQ+6Dm/PpmmG0hVfm7zRqRZS9ukxQ5H/nrtSJzqWMdkW1KXbrq3fhJ2gT1bWbl37DECLfED8H
DvQ+ZQdOp8lzdW2Vv2ysZrCVH0vHla5j0sBzsHn+gKLSZ5BesAfst97swnAIItg5e0+O+3iQsVoe
Bob0n4NIIVwx2RFkG1vWKqdqiKNFVd/PCqWIR5u9yLh6OiyrHDA6DlUWQITsj7FpnTMO/kJNyLUR
FKSetqHRVZ2TsElg0s2An9+Urq13rPN5drJ0vQKu7ps41l3OvuV2JZdrVAQFUpLAO4ngzdNqHUjk
TSIMPEQb5ucVPT+ltgAmF7F0dokI0z8mMzAbgqiqYIv57LgsTvKXu9hE8C8fv1xoNRPtUZEkUovz
k21g+RmXePx+eyaIV/+ex37XEs7omvw7f77dSkJE37s3fWmHs7nEWtu+xFXPX80fjkL+x9MOqui+
FGYYGJSocSzaSNgw115KhtTaXAFKPg031WevCS7nvk6b1d6J9LjTDC4kwk1zFyum/iz2oHwVELSw
BXTN7TW+kcuVtUfmMWJA5VVX6J3v535aYrOAzqWh0/tri7hwrZuNByJJOZJ6W0y1+ChML+4WsfuL
wwsQgDiJMXZwxrrbqCIDmF76a17Woe9mfQ6fnmMrlteJX+EWPk5KDynGD4h+92vA5s369c9zmEmV
dYLd0d9H6iHEar6dAimA+IMEeOfVs28Yhn7yV0LIIy1eFK91I7vqxMZRKe9yBikGTh/23rtUPDNt
jWcnKQdfhlvjySzX9kDlHKe28u0cfcfVbGSkvlUKmhLNIcIzRwkIwTc2GRtPVcwG2lIPoPKWCRdx
FfnKCJk7Ntn2lKV7I318q+XUBeT35RsgUSJk6dqHg9cVFAaMhk3TMPf1uvOZgVPLpTkpVHwsMEbT
x+USNcZpxjLIhoBiChn7jNCOLR9dDzDgOgxTz65i+e0y3llV+PyaosPeTk5fyTF+2M4u2XOOIz7G
Nt/gKMXJ54S16+Ib5e9IBcfhlsYiHKOELkkv2uvT/RRXnWuAwPRYCMk+kkHFCqzNV5BayHEhIci0
sDytDxQDY7yO1Djh3KyvRVdWipX33+OathdX/DcxmT+pZ4jSpSm3kKbQ2T9FQ32Qdjlp+pTlryKr
kh79dit4SFc2mBYeX6x4Chm7bp6a4g1JRj3Fy4Kb2pdMcvcPyCWgxB4asAK12xacCxQ7XailSMLe
oi/b7wakrmtzZ13QMAgGOAjtb8C/mZqvLabRi8NraDT/8iUD+0XH+S/sTbOglgO2odmt1MOe+bXe
swRUJmK8RbHp322A2rExq5zBrLRkMWVTcSLW3gkwLmmL34Tjk2qXneqMf89EFn367GtoSODs8weU
6NVZJOlX83Q6/W3lUgxEkFt4V5cjsihwPIP9w/VVnywBSypEMoUhmdbmGLq9S8JyUiYu1d3kIsLf
EqfB6aqvDPnSxT2MbgGaYDQ7sg2RHEMMvkBW4vDHQe0BZKPFo51Dt8Gvilw4lT5J4jQcicekMWXi
FUkrI/lRnsLlMmpfqEeX1BApRIp+zFtyjbbHvTp9YfNQbavKz2u6vd1JcRXjQPvCMUoX73nWsbUn
CmWdj8HnYgdKZf/hyaqBD50Llq79hUnXhc+KE9UVK+in2RsLrG7ZTxnCULnrd5vY/HIAA/FnTp3P
x8FPZfM+Z7eEtZOeGpOges9WxIr+OK6dbO/fGznK4W/6FXL6IbcCOYTFQKaLKUzxFUKDK0U6niNS
vaXvBSdyQwsLeu2gyeWN+hcNg4Jw4zwgExeRYiZmiQzTuw3rfIbbKbnZavk/y8bc8PG87rvvZ1N3
mVQdF55gGzRxztR+9m3qsQ/gOVG7vPRMfwvGetTnR8gyC1sqYWPiG/qWuMUyhk5F5WvD5uxmNagL
T9bdunza42/zT3+I5l2sfjOPXKb/sxF4QTUH7oGujc7sKQCjGBuZ3eYn2dn9HP+7uhWjshaFum+1
JTXMEfX+tzmtQg9dlhUkDE5KIltOHwPyT/QPhjI6o61x75/99QJ+MBq8Xkfiv8EF2UMp4cOj4ZL0
2JIV2QdvL4P03DvrwFOYmmLv7IYL86Mq2u800hcGA5TCt01i5/L0+uUDfDw/P2QfMzDsOmN7Hn+j
vPXg8cpNpoOBLU9bXwoLnVIY8wg7EJUrncyfVtYBJjVpY4i3peHihN1+STUy6kF5zgpS4AVrej/C
9hEK6nT8GGzbp5+vUcGAq2jzOrnEGzKs9nZtwIuYAfmKztOk+lBqFB/PTVXkWr3g63n3WUkSNd3i
XutrFl0oLJ9eVZGcyp3nsq7L2xCExAR2MTCHi4lZ7BjTy1URU9x0nPb0pukFIti9tSmPa7v67GLr
hMdjiyFfOKHoqqjA0GXD1467JTPqwb36oEymmv7rraoqVZqH6Xc5XRd1Nahkp8RYyteEbM2ETvOw
CmGEYgCFFqHDTi6id5fwUpyXDWAAnjDpT1ywR1hFyjRzpO0UUgOkubBgz3SpZVTNw5KQbtuet58v
dCOewmgvJjnPN+4FPvJoejzCN4rzoEasDUVWHFDHfI5+rhvwo/I0A4lLKqIZDi4MmygYDV2woSM8
cNVsl4LX9Wy+Ek/v+t0CffaJN3IOQV2AKGC6QKP0l7veMcjblml1nSc1OtQ0VWsCleFyrf3RkJuc
V/zY5uk2KqTwN7Q2aRNer3HUNE3wALx92a29ydFRsMHqQiL50zPfp2ZaRCJpQ4Ka5zLag4XER4kQ
ZV3RLfrx29w6CS3aV7zYjBfp826CUPh5CnedYMVofoHIgYGLUZH+qqBcHb4ZEfj6uuubXqCTnMAG
T4XlgwCFsUyuehoMeMVR8W+vhLoSYuvHFYs52+dvyGja6v9vNBn0LyrFrb3fBDvAOXHuiSsBjaG0
kDRYP/DkkImkA1ObL0wQYP5IAKn7Pg4ALxVnCXFWvslSwWdYBgYBYUuIsWtDkFZ8ClNhKOjsIsED
TonTkUF8ijQgDMk9h51ytyJhFF7AfHPotmLxOGb+6Uz4Z6hfuq6kPoPbqrK5Vd+9qDF47lkmjroY
O0FCrjV4S+RDzQh1DZ+iLWoIpjGxSwXFj7hFBJ/vB9CsgdlPV3Aktir4a9SPLGhv6+CzwWH/RIjL
nYpIzRhVC65iflPMBvAx2Bptkljbi6aexaTqaDcE/LIy3bqmiaMrJa4S9zk1px0yTBtLrO+hA8Ek
1tnrI4X4fK+jRp3WpIXUyxGoaCygdka9al776Z+p5jOCJTb0f/AknJxSltlBAv+rISyH3m6Om44o
MNGNzEQS9Z1uJX7FmpK5SnaFO8Q8h6u7aFsxbhvxhYGEySsd8dALlvbd7lwPx1KDUOhVIk4tTZDx
y/onWixxTEa7a31OZ03oO2z8MwGoqUBuJ8U9Wd5zMAWFLer8mMEmxXveSOEfBze+Xtq3wXVGCW5+
5tmbk+T0RhZhJl14a6kIJpYfzyiEbgRXxPL6kAE8e2RjnJv1/GvlSiSHb+aEGw0C1FRvsJVmdWOj
ow4oDktEe/ZaAE6scDG96/YwPFWF3h2h9GUZpsmTf4HeZmwBikpZ3Sm3jQy73eDtjYMcYdK0H4I9
iAeoQv1EXcS/uIoe9CUgag4ggsYOSgXmjf25v+EMYIaumN0hHTVX0tGJWXA+QinP2HMe49fdjSsH
3huIuWbp7/H7ytd8RRlgAmYjI/p4Hz5ETsNBj9mOB4DVHn++vH9yooXs7W+7/J5q9mwXXyDYmU+/
+cT8RO81fRzZ5aMr+hGe5Ha3zB+J1sQ2jnAEXEsWbsozkL+PzN6EErr53R8o34NajyckRIWt1fL7
UJRgF8f7QRKV1Zr9mDx6Coclwe3Kz7e9xr+9HzZO2hNWC+mEBnO6CdmUU3WgahwZOIpK66NTJBBo
ddas9ciu8zGt4RfPS/UlPUitiiNheE9tSL+7I084uXvJsJPem/zOjgS138tMBrJnWzc2mZ2vucTv
2UVHWuEo3a04wCpqsSfn9QK99ZRxfucFdmODGVy1Er+jxcSPfXcU6C6tYwro/Pa372pUCCycHjUh
LWZ1G+EBw4zq0z9yn848DIRBEtq5N5vX1UgCJsHZorAkjPwexelRLA0p5zaNLQ84uDklEOqbdaNh
Futb4WLfNvnaX1GxUVPVBOUd93nXZWQwjE1yVaTZrJPuRN0A0oaLlpph8j2yk/BxscRGuF9F9WXe
4HAhwyOyE1vBVEoG1qfezThp4Sxr9sB9jyPKsvrBoDl1asJ5qEW9pCKHm/mJSxXmK8WqDx/9Xlhs
/MychnLbpYQfPTWlJbHCGOvc3Ze0J9Dk2Yhdnyr7VoYkiDqrrL22Z9uhbX0GQi1yWM1/CUTuVPtt
2vm938xwAgWHRbfaTGavIU5QKkH0b9cPIlQxE1d2WU+D8n5Dn7XZMdLpH0TcqKxUxe4f4FeKVcVx
GaFai3+VzgOiIm4rLA6vzDaiuP0znHcJW/FmA+1YmZf202a5+EhAQ1DPfCUkrUUxVzZUbYfQwn6O
jLtgz7E7Bu51m2muRRWxghg9ewaHjaK6umn3KxbK+Es5mgq9TSRGcLiZar8D2COGKGFb8EowNYKS
r3iUGGtR7QoTyZy911pgkVp/rC3vTDghbfBb3oFmfc8B5Zp2vfWXmjMAxz3vzY9islB7fZIny3iJ
NboMU8INaTeR3YIT6Gul2KS6zUJxKGszohXD1KnazbwpVfYTPGTn4g3MlQy0P2aMZs592wf3qjxK
V+ljF91ZIikPDykjNx4RUwUqLdd6Rssxm/VDwYlkI5RQNlKMxnn0GPRqXZ8+9ELEo9qpL+qlAKt9
iX3aOM7FmANYseVwKFyIlqpTzSxA8GuSmsWtb2tt/cZYmRjZ2l7cyQP4hxNs1J7/J/x/WvCt+HRp
9Lt1FQmllDRvIJLtMQFNTD75Bnxhaa+NzpZi/UzhZC/yt2tEY1YjhNkpT2T4FMZGALGYVqVFweGd
CzBij0/fzIXt1Tqb3vOxHwQ6TQaAo3VSlaYzREw+qXSB8Cc0ZHa2Ax38ppm+FCDBvbfXVQNhqHKA
nBxYrejougpxiKWl2gC7Q8UK0JmfUpvDM/vm6InXYhv67DnrRgt7s/pffdCTDQeRKrhlAOr/97w7
oEUEBGysjh2Q7H5sHHq0KcsoGfgyzrE67CMZKW5+CUOQg9wNAF2v/bWyODe6iuqALqF8efCPeaXJ
lg6aHhb+spj8qZO1SAnJRm9Zsmackqh5T8Mfxx1h81fohYl6o96vMRqy8S4gIcUeN38U0fqYsvmW
FZAO8Q1cZNnpPVpBgdDEChU5jbZ0uMCELDCCohJkXR6knA+x1nZ9KY0MEL9WNG+eK4hQpRGxywSR
u7euyUlLaDi6fULtJMGrX9+rtqrbkJB3XSlDaDlwkhbncHlWx1Kmxs5tp/cOVwoMebnASn36T2SI
9P+Ym6RlZVAeuYdEaaJVbOaoV44FjFGKJxUDE4mdj7ZL/wFJTFF73bQZQt04CtB8KY+/QhPrGM2m
6YXrW6z2raUpYOAU6WAix9L3f33iiy024pxHMg/GjaL+4yItKGmlcx8lIt2T4uJLhEsJfE0GWgnO
Ag+UsPp3GnQo99ch2NuyVHSP827MUI67m1DKFMEiyj8H1kbIxS3OzzY8QSkW5KwVr/FvwCkLnQL5
enJgygeBjWLv6ulR9tHaD8GLQJaliKuR3bCUM/ogaCneErUpZvlik252KCu6RcGIt7bp47DJaoFV
CD+j4HHoAfK1sfOjGFJhacVB/N0/ZN15ksLNSsE98smn/IBlXu5vDr7yZut7F8r+96kRBPp73Hql
hFMndjIy2LRSLemnrCZBHvBK1bzf2lEevNPQEsMTo/5B7ClR+eGDnc/b7QM7YC+Ljo2mT1d8JhO8
cpyzHcWN0Yfcus+0FoBH/x9F+hE9Qoi+Nn0AeY941mAAaZNEqlJOzb4NqB853q1mwiPn5aSCoWce
wD2D40UlmwXdwHJPlsiyzPdT2OnZQnjnYTkcCYvvhQIkTJU5m1JkCwxiINbdV1M//9pL9ROco/zP
OZFi5VFObYpyQPJpSuPs1Q75lOrEChsbKs5CtVYVQmTxnZdtf6B559N/EetCRqyl/mHTDH0CYk3s
iLIy4qSxgvu5P/HDf8cjfBLy+OO1KU9QHU+emHr6K4mnI6+sW6MJ9PMOdct69XcwzzBO16FhwNG6
UxPFwgq4FqIxwvmTgHpK0vzSTn5xAyNE67uVSOjGHPZMfceAiJtUYSNX18QNvpIZ01z3QdpXXnYf
Bwklr4XVdozdoZ9/AQxDBbL5W1WLTq2+vXvC8mn0OWgGLjN5vr4Dopw7Rn4kqSzNc1yeTshI7eew
DN5aXhGWxsaknCexytzI/8beuih64TtayMmkMpHZ4SfKYqkaD15DsrJYO92cXnYNn+z5kxW7XeLw
AdkjQY8SVrG1ZKU/BwTEeIlLa6aGZNsJ3oz8/ED/ciKF0eI53YtzjRBKoJ0jQ8oisWWV+CwJtyFa
S/DyQOlp5WZMdFaEF0wFdgnztRU5eoQSO1nb4K+JNfHHrs6TCRkKJzJuRlZnGIIlvQWy6u6vi6dB
nk6KXRgk5yUw4Wk608cyqB5N28d2zERQwUshdCoPA3fEC+iNwA1akNNn92GyHnvOf9XFFXQa1St/
o1QurOHbZoWTnmqQ48vE0DNH/yymqrt/ZsiJRlv1f/PzGhg3V9NRO5yxEtNKYOi4E9x7Tln1ugOU
/NlzMecbx1YqKrKF0eE4UeCRVyVuOOm7tU73h7hTTL++livvXBRcZ9Vw72VDw/UZRwWSqToS2GFk
/5gJlTd8DGKpa9hcbwMNfAYX7qRI8tJXhFjaPoK5fjv/qWrE8WIwGxCdhRUlUjzQULZc18zPKKtV
KUXim8r1dr5zD4AUZCprZG+ARJspKq0YMiVmYbNDHoASa+lKaXD5YEOE+ura5A2gaJAE4TliC9cu
7rBz+9v6vwsixE1u8EiRqymxnwvbP4C50AcufQfUJ+h9n3OVhBpRxJU56fJGh/iBysY3fMMKW3cG
jtu542lXiaTCC+BACqDpVbLudsZrVzhDhzVrrzk4qfkfWNo8q9pZIEbquHoN1yAhSeQsiQp8BafS
86JX4wBxdFes16O/vXO+BWOO1H1VQU+iFfF5g5+1agTrhxwWFH8TTpg8M0hb7WX6Lb14xqaZMoFI
2CSYTHtd2mNXjNKnHniLzRbmVKKVwRcE5G4cr7fcutHv4yxQXvn0lqaxjfGhbbAOmwf7j5ZOFQJp
WNhfoDbXFIo73OHBcJ1JOWhVw/Ad0u/xkgl4RXLoWm5p5pKEo0u47F5LG8vC5CfU25zNQCcUAbQ4
TePwOQuTtxWTt8GYm/fGHg7pqzcfcsr1nMai9jFr49TVsfpw6fpBEk6eF1JAHIRUDq0SSe0dnYaU
906Zo4V2sYFQIp9IKOiDkrNvO6tefxUCmrw07t4zFDlpYTzUGWJyElAta+GgyHVu5Csg/iYzpwhA
AJ0OdAl4Jxs/7ksE7k1tMhDQXhAcJKK11Y8/wpF4AwyJQK+ExueBy4lsicPZ63dCIK7Vctg8P3Ex
uK/EKNCA9yi3f3OxsHCaWOFgcA6y2m7p8ysR1D9oUVzRrDtI/y4Xix/NQyvXKs/o/y2IVKwURF3W
VDt3xMzb3BV+DsXpHuM6HoiLqHWq5VaGqQmU3L2pl63G8vQjvn71n2qsQ797uWatRKclg91tNeeA
lb2GEx4sqPIh+c2K4w7LyMXnQLw25EhpgQsBwZ7aS6LLccVQHPR2iWFEoLUz6MG65vxqtPH9ZCjm
8WUCLdsZKylvIWxH74/7yRSx93sWfRwLH2NJQpQRNJdt83aElrlEDtBPT6IYArY74Sl2CDKomNC3
4pBIhiZY1/LzgtSzpx1UREQrZ3VNLdeuHBqAU7CdtILQAsUSr42AByIxQnuf3pqtGGM4P3WNFu0L
79EeR03/nOleVO6VYJ1J8TmpvQWY1FZIipmI7alIX/raCNTlkk2IKNdbgoehI2T7JONo4Ihw0jXt
0Bw3CS42RUXWZXeFaAEwtBhUYIu8ChU9FBdpZztwDiqcRHEtKtySl3jLjdCRkBDFqjeQXlZ4tTze
znb1XjakCKygcMqPTQlG8HTefSPr7KZUwUhMJJFpV8QSJhrgJyoPgo+OlxdEv3ILmGTt6TusGSjD
xGc3MWcADry5ylta6wlpTeG3RGk2R39dTYn/PQSve00xjNo/RcZLOkoiSnK63cE/hJGsAdqpLKY4
t/Kla2DdZAee+hYZvpRltoSfj71HCv0qjXlFM4BnxWVvrkYPF2HPSDj7clf5J0yE1HeSNoP471fU
+fZLrdY6JSMgSfHBtB0X+Hz4uGSCF2KPXpvV8Rw//dJwdNeLAlc4YAltpANpMm92OwZcrB25wl+r
qVLSULp9soX54L6mGwEi75I1A4c+vS2aha+MsAjN+6XDj/ncasr0V061Amd43WUg4Y9D2HDVnjDz
qpiw6mqAmvBml9ISv1zXXluWhSAUETDoXdbh67F1ja3Ht6+Q3hmfDXnd6UbaX107RwRYgtEnYDA+
yRIxzK+zeX9Rnmr3P5+RG0i2PXNUeEKqHXrFRWHIlwtPRQ1V7LnPBGr3WDGSmaycyLzi/NVlxo0Z
jIjqXs9pdkFobTwSdRc4u+nUXUhkN8rMGP0cJKyl3egHJ3GvjOutjur/4J8DUGEZYKizGZ1p/zs2
ShnfmSvNqDZ/xkngFqL9kzdAQujraM4/rS1tgX4jJq81fJnylaXEVKyP2znKrGAXq0i6xU2RRdLr
vpcW3qx+zo26jCrXds0xQT9srz+VkQqzZeh0nmTTsJvq020G1GDlIow/IOfVP0fBZFKAevmTy4IC
/pUtYoAOWBPm3UJ7SxdRS0gvZLdQdvo8QFt4c3VW9W++CUSullyWne6765m/7U6a5bNWOMF6g/61
EgYDEPN2YeQdWZ+8wAY5/+USlYc0vjvK7xUUKjiKdNXqXLPmIGH2mTI9CF6rUta2ihIUsg2YM8tz
x+8uV9x+yQoaCEmyMN7YKs1Ea3MYqaeF5R0VvchSIbOSwOixMGRxMBDvG2KjhwDiK6nSjGVSBAqW
VsgM7gJJApG7odpFO7GruyOGP3v69SiKYGheMaHen493K1aKQZp67KIVOynjgRwt3WygdV1PSd/7
l0IwNLfpKhfOQRD+msVVSfOJ1IeGGVzgFTkULCMOes5gET6ABF9SUrjSqGsd9EMJraEg4Q/3j+DE
nqyKJdy9J6F0gAiVECrYD6rbP6fKGopw4jBfHnYSRtnRGPdMYOt3MkfdeqtXBu0R2OiLSsKXkr4r
ERgqB8l24R53HxrSVXJ+teRl4XNNBpYMX05vZ9SBOzOBEn1AyCaXNL7W8q9ACWq6FcMo+H1ro6gj
Bre/ftrtvyuDIwdGgkhLvz0/C5qWPyP/PzN1fGEOvHCIV0E+35i1NHNH3MLKMI5ausBTb04ak8BX
7sE04ahzCVGEFeq5bDjdwpBPIKjRKS0H7OkD/MxpP3soyLkemeyRdC3NL295XfnFTBrdHD5HOmBR
zK3mas4Ppi+l7fAmfRmvAVicoxqjFyV4IItfu2SlL/U/6L9cmTD9bUDhwj+M0Ruu0/Tjj3X5KIWm
1e2+qEjrEQpzLOzMWx1nTwBntbuTmYWX1ELpTSOt45xE3Tf9o1OHFivibjD0it+JCoBpdrLu1aL8
Lu7Pi7v+RMhwd8EYWCwSxn8jfBqpj3HVdA73YxzpJf62qdY5yVCvOZQERJScj7QM1zPtL8aMXpFS
BlAwYagyegfuiRADmO5VlPuxlE4hG1DJ5PZ3AJEG2cEZv4EKQhRn4MIELEa6ZTnBn4UNI2DYxqvY
12GnxNxmwO3QOveOQjSXNDCiWBYcGuZiHweDDEBlfkgk3C6+1F2Iznwc0j9FLMmqxrm+Xzy5dp0S
6dW5F+6b5od2v2JfxyMsGNnQnAFB99U2pgSSLPdtt83wOFkx6ememAMC87StgQVTJcygcHIS2AXs
PtxmrA02CIV4zxoY9DWg02tJQZydRNmHin5khU+m2t8V/SZPRYJWqv+kKhNoMz3rnN7+kZgBbLZK
UTdyQEoHyGu39qiJQo6VQd9GMBoQIGA0OKNsEza0TIhpmpEuSwzo7RKGicw1ohqEDOhQxEMr09fx
6kNKAA4MA9QvNz9baFnNIu5Ig7f2L68XXkFkJrIywwTPo/QLTVAz+cT99rxesqEbsi8Lhb6VE/oY
8sytKW+emTDrZxKXEt96H+Ot8R3PwJvkshRcQLIkumj2JiBLsuk/MnM/UrI34dq8HxbqcyMAN4Bg
01oScvw3huoWWwZVBb8xF6GCDfmd9mU0iiWZJmX7iqiWH+XkPlmUsXk3FIDZzCnZnx87MFUNn4dE
qypuBVuAQqMvO/He1mRhD1qnu0r4TBQLiT0duWS/Y4yv8IVB9aHnVVIoKu1b86TRUtSUihmQ9x77
x/tfUeqOt09dtOr1sGcNSx4JND7u9TaVEW/pzHqmwfZVk52vwx3A2fT+l/S9odZlHfvImEnP6zDr
WYl31T5PHcUjfnZ/uQ08F17DyfmUFJ/Yx/qCrH732NeOsnmNsia2Y75pR5LmxEhFS7qvf3QXZDNl
6JZLwhmWfi5JCMH/szRTLfnrBaQl5Ohexxw9M+EW8gzD/ecjEy72rlgIFFxrvl4D78OeNks1q8dP
x5JLOOHCssshWqWSxp4kIS+rMF19k8mQ1j1kCwcgYwr52AGNvKdkB7z4hvw5e/tS48E5og2Fkz48
ET7fd6kCEImG8yMVNIcC1KLX33c4yITjSG+eHGXontmkkC3q4NnMNoo3EJZ9fiGlWtAxKIoGFxHF
ZGfeHKwpX5b4kNhcIj/5nrXLRmMHlg+SSIzCmSJQDfaFnxv3jvbg3N4rTJmg+WG1hDRIrHNYzzl3
JxfteD5gnY6odZzYBMR8avpn3H3v7CuDzL6dbXSKyVZt0oNqz39RYJPW0OLS56bK1iOcoPVbiprG
h0y1s8a550GKPgvfbYkbO5xtRWVacg2XhVeTXgWzUQcEZVLqzJi6OWTt8kKFiUfW7XAI2Xpx42nw
b78AKspkNss8Boyz8dT5+sjEkG0yVGvJfv2VDymWayW1xi7d9i/b7i3nddH8kYuxADfwlQVYdZeb
Pm3/Gb7Bkgxg9i4H0RqpWsOUloEEOOFv2aNVnsTIFswOd8JsyayYT9TCMM6vGNxHqGmHVKG89HE/
7b1I/6VbwHMZcbwdeW34ZVwdYIeHz7/F6ottKvM8RV6Ia7hVc4O1wJWyhtSZDSM2jzW5REeWQ7Og
b70OqruyZ21xD2s0u8WlYiopZ4h5k3ClfmHukgItumQl6GdBHBcg4c1UeMqFF6E6+6XCysyzgNRo
ay4zC74PsO/ipEvTO14BGn9Py6Zc5/5NfqeUJjqA64G/QMTAO8Rn4nU8xQ//9LG5HFX5OeMbfbWV
rKsfnPc2zPkWe2ot6gMuE4Nmn7YhKO9ErI/JHZBDaFrjutCo3zGmUFhV7jKfWDBpzNl6fal3l2Ba
JIGtapHoIYUTd4LwKk9WeqU5z+VHTVZqYac33AmsqNClkbdkcm+mP3zQJg0/U9NrgiL2LTWDkkXQ
p8zOK/BVq090x487jOtvBO7hybRpd1yo43TX2FEoyl3OK9qEX2yTkypNoAZGf/zEec+PVwgLlNAv
lPP093jEGwxlGHrPTgnG9hpAWpVV2pmLKkcmPb26lDRne+KICk1ZMTQSXal5DeDv1DGs0KKrNOeg
M2ltc5nmUv420xXzNXMsh4C6TVKHiQzP8u2mIo0JLoDJCbtymbNRZJVUXO4EpbsePi2kO2KD2HrB
8a1zSGZf19+uX0OhpsakKDZe86sKhI25kper2dDyNpw0ySgv+L9P8hXrbAABhieehCmXXMZQ1acU
v8ZhgDRPRfJJbEwdUP/expBP4wOfCTyqpRaa1jB3uI/Jwc3bSthZjk9RPdu69k5MyOW3aK1RUBDW
VP/9yW6i6kMIjMAPUywnn75lA2CcAM24ePytSqeEBDtf8mMLUptAMU9+KlWE0qoi1cbrknmBwk9h
0jY44V+UTePXVpk+8P8yku9X0M+Hhmr2cz6UsynYlUlPI33zQYmsA+WTk9UbO7FaYxSGTOyspLoV
Cb+ql3oAHfz/jII+SI4YEISK8/44qAPhhNayQ9ICOmrIbBEDnmoqe2Bf79q1mbkSUyR538XBSsr9
YFD+itU0bIZDCRtzX1mfaN5zXgwrEQdqHyqm3MGnqmrTEg66bjQhD2LoYKwoyigX4RPHbP7BXxoI
pmVrcQkva8rRSZS6x9mnDEa/MbqS6M2NApyjS5O+HFC8qE7Wzvk0BrZKsF/Fl90xV5uPZV6koRFD
CB4iSkkNwifknJgKSPpGyG4/6JbaQUYJ9O+6lL0luWa24EdXpUGVMvdUnFmNwdUv/C2GRRzhHj9w
LYU/0klYIZuoZ8ZIognvb8E+kdE942qyOQ8EtnPSaYJqI68+31EkQkAz+fbROPZylY03c5+tpIkm
MUSvf2PTdj5DVoJglYnJr48/CUKvzyY7iQoC0sWLOWzF3HoXj6NodgAEbTz2r80Nc3TnK75yJuE2
OZ7X21XJ74SnNYPtCleBHqpy6gk10K/DXXbIK/rPkSL0tlTCGL2AL4gjU8FFClc3d0l7IAj9KSpU
iRzsAukIF+Yjm6AOPqwZoVhCrWKG6HDKVRX/FwmsYnRwtJjxSZ57FpOXRJDrpS31QCozEIIowmwy
cUFISAI6gUoJJrd9YpqgsNMlfpxy3/JNjKHjuL3Pely09YRwXkQb21lrdfaAoEApxIe9lqK4EBpp
yb+pfUk6TjlT1x1dXAUqpoOLmLAs+pkN4kXCgFi5ZQPyHQQt58yy1ZjYo/12eYPNORDu6dRKMosB
xJlwYfw0LzNtNFMvj3jVVhWYNHpGR7fjEaHqVTS60+oqVHc9cxIJLX2ZEWBX0236I7w9VH49DDtr
8nTLppX2lu/Mw/SXqUlv9O8Z0BbBBBML3K1CobIZZT1fRiikVnR6kRJXNrXfNCBfvrs0pvCmKUy7
l6HQj8ZrWPUz4AWRmoZFuZvBNyM5zqiRlPshVz9phsWce0A/8xI1vx9MYQZfhUSkT+xumpCza/MP
2mCuMUKWLpo7TZ83/CHl5UrwAtG2uA2IHOVQqX78+NbJgVQyI17MdbFqwD0Wb+WY+iPOPBbhgpwL
8rU49Bcv+eGUY7LzV/Sbn8TAAZTaBMGKipShhN9aiii0a6e3ffDNcSVvHD8ySHO9oam8Zuh+Xh3d
RAyHjxrdQ7R2+cU9cy6xdABa6ZMm5B0oo69/jux9ar1sqMhysFS9x5CjBnLrxDgrPCBo3hAFVcxw
OJgn/8HW9J5djAMRnaVjZ7vz9NKaD4xrHs4F4E6SIWkYYVfSVxKO9SXkCuZlXrLEQhrfo0xUYmX5
OQUwzfWL+M7N4F7DAZM1G0tK/t7qaNKw0wrmoHlZKSK2mdam6BCylsB0sQpXdVvCsqw5230UsrER
kNw8TWXgHwvNxFudKH5hlBHjABoajsgjVshpidYQ6sTdub7yYyEspJArD1vyfBqM9EmjvjUtVtWQ
XNOuroEo+HzgkxsoFTawGH7+cPDrcT0hAvPG6QvddjNZNRPrU+TzBEbANRm3utacqW4PZRbLMD7S
DH96impmwusVsSlKvTrSxVUIZrRWl9eZ6gVRV4jAm8/L8hbXu1yECj9yHJWdLWPBFwbwe72tj8ja
nMCJb3Barphn4pi87eBwj04w5UOgMimP7V3+9VBUnH87darY8ck2VSTyBC+fb3TAytEt1nWrxdUz
1d8cLh33wt7mpmN7y2KEm1nZvoUUri1leo7/GJJBcGksg1T6ZUN0YPB/q+/p3pwAbQgan+sYAkqB
8QQUGJgfIDU+2S0f68gIWyvGlbM35SCeygdpMX8ltGBMB/uW7zcDI+5BnMNkANRltKkGJkJT/iOQ
3X9k6rE9hD3rqQnXqrcz+eg9kmNSV+6JkpwaJTl0teJBg+Bcmb591q5ClHY+dCYncc4lVqRb9PpV
MF+CoxNvtut2ym190vUeG2bpA4oL4chwVFUqyVYtEsiaJJ5JYXgvnpjqzkAUGqdVzLX8JfKia1HP
s0yV4JL/ag5NxDPs1b3NhY6biGW66YtB60/l80GpMaXHV3UX/IZf8WxuczyLPlfmeH7bvJ1nHvGY
IX0L3qUrrTZ4FIhiFJJLVhaPgHnQS1qGyJ+fzjnX7ulcZOiH7GQf/wrKuz/vmKmWZrdgzAnueAEN
f1D7P5sBS4gcBdGdwX0LTSxTfuSSpDbykqd0cbMPzsXpx1tkRVxsKOpVayKvMJkJ6TbT1PRi299B
A/7JDvQVB1JhnIMH7GuqORQdaRc+ac47mXgYG6CrhHp44lkCdtgra94DkCjkF2IqbHbSDtQQYFaQ
XngaYB6BlwNKE8lnEcnLh2zHwo5A/8t7EzgphWG4UtkJIwOJMiMimD86JD9IQn1mvoSZpCbgdPdF
o/UJ8EDRz24phG/+gOW8KAtIoLQf5V+tKwZhDITiPvX8lvSGYeS0o7jiUBFLenmB3Nm5yPxEqF87
IQ3kja3WaDUpo9d7l3CnrlsX2F+mpuAGaVq5GM8lYmFb5RsWSxp7i3+Z8G0D5j1PxIcwZOeNgGtM
tbNqLb4SK3IzBOjLWcGZtEArfipc2im9lRZgRiQl02qTPk+Sf4EixzGEMEFjTBFbda+FwkxikFL2
0BJ0K6kDsgNeG7c9KzohGL1pD8ozHbbnePxt77CiLs4P7Po0pUNYV0zNGtRWl+ADzHQMypfOuHs/
DDEMVkYbtONNBsiLc+PMaaj1RfrEnexO8jcIldrSwQvTZXfqy3rQi8atIO9LewGP8/KUiiN8kmuQ
+RPb62FMk63/Ys7kXDkhFAo9hkMcUvBS9hCm1XNeqfUKQ++iMVk6cclzV8VBYNk8G4F6qdJhbkbT
yd2LU+LWpk2vYDsNUFmZeRc4audnEZbqnqp57IQIIE9hr1NbkBqOG1lBdFNcTSpWTNTJCp31c7c/
WrrO4zUqbqxQcl+QzQhOYC6WQT//80Gz3AZPIWKi3FK37J88EIvtY4xWNSKsD2eeCMyfNQCQwauh
75jutmqZNLgI9rpZvN1AB2av5jJN9spl8GS5qWiHpTImleVgKPkuZ+Um/T7y7PMLvAACx6Vhaqs2
tF+j5+LRfz7CsFCJD33HzPjvC4W8ZsftFKIoCVPNp+wnxQzLNeC4ropTkZoiTF1CxHndWUDzO4vS
rtXUM+AP6P13ljAdqUpUeoGSqXiokzVe0IHdDqrz6bbbXcCTXZfKlSKuxlyD03UV8s6lKeJNAdx3
V0gbjIkWmltzGah8htQgnSog80qIwjlAlqx+4jWZArT+e7bjU6B3xtL3bNyCtsSD1TBUAXeh/KZi
Ks0t81L+xkYoIw9+goU7Q5ZB0kAaJzuLbC61AWoJFon2Uq6yuwFPdd+djRzyTDoPFMsoAPr25Z8W
XGzEa2DeNgJPasBl5EFNAkY7vWjiU3oGSFd+3y8SI6ynM6C3sAHLTC8aTmwC+KaORE3DSAMEAPw9
LnGBPODAGMouIkgQqEXB2bTGLKOO6Uc5qFHwn8Ae0ZXv0WizevC72uWhT5uE3TI+dlxIsV0YncoA
8Dp9q5PXSWXJzkmEF7xEZEeUP7x3YWSggqsajyrmryN5CY1cOdk+vhowv0e0+dSg5csLkeUkTV0E
CYfVsBdbeInnoNO4LvPLoEPr6PQQUK9FqfbKIiRwC8Ae4g+FXWQAMaJb1SbZcAfgG0JBKIfyr+8b
MhY2ZI2pg9rXcygYbcexfxfCAArQzTuzsO4cXWkWBw+Qe/m49V3Jsi5ii5MzzL3L2BT+ck1vbcDo
XzSn5FMaX/TGpM+S5D3pdd2oY4SxFNpF4axx7hxkHOnZLhV+YvQLdRBDyUmT0MRYGRN5mNViUYtJ
ix6YkiGVx8cKzoJ8qvom0/XMqeS3W+cv9I0YtxKZDNPvlkUrL5jfPtZkcDB/CUZ3jfczBb93nPbJ
zOWdzeWxM6Q29AghbKeQkXbn6Iy3FizZ30s/liOVjr0BjZ6TIglBox1HXHdeZpkqsDIfvlRpl/sE
ycQLHpelj5pLr3hQczSAfhObD6migHPyLVSvwLJemCAstWyTRsa+l5qZEatO2IiDN2Rc0TgvL+mQ
wWsCOQq38VnewnTcUaFNOa42xCIX8SvnBrtYawSs/RzQ8WgJIGFKV320ErkKuca8//knHv/0xwd+
Kp0BCqmnXjs0P4x7xTxY0QGQS8eu6Wbnv4qkA258oawdRyP1fNvm5xWQmD1f2QXFlf1atYy9ftDc
tiVOoRuRl6gixSzFEBBm1gUrYqrFEeo29qNsd4crGuOsi8ikAfDIBSBunnWujkIjvNfqGGHYDoyI
Y/h7Y8azTzITH2LWZfOzT5qBuZuC5TAhox2DIAhg/gOzpO39BCjZUC0F/MpThojMC0/pe0yMjBTA
q6mjGtkumd8o5ndD/u2hDjTZxz0GD62ml9RoQThE5u8ZEfjwpkpEms2OhkhvKaegJeQMUoLb+vTQ
0IUWKV/iovG2J9IyXBFadX2KMnEyxpxw9rsp68+4mu7lJR88CuWJQA+GmCSDUoXkmEH8g2nLLTW7
lAX5VB3+EUaHDYkwFlp8xHDwdtnwQo3d5jN7EkLnlaAD2NZEYglgMWViobAfPX2UCoFpXoSCKpmJ
a6+LZqBRNj2QsMkiUnPZjsCFxNKMqt3HYSa87OW4wxdGkKDsnQssBhGrnYUaaCxl1ssSZX0sqhev
wws06fwkAuKu8FhTmTpkM1CmuFFw9uc62qy4rUdEnNtbvpauqPqY+P+qFxzoSYLi8aeA+ho8jRSU
A95/gwwqdgnYEZ9oM60rxwATe3LS9l1cEAC3T8qsW8JPsUbYLSaZdRk0HOJZDB56kJefy9lmiHIT
j6qwWcCKmBTs7g7a6p3TyAeqHEk4GmLvS5qXVc5Ad/a9GPIQCkBKPEmrDorzp98SIC5Rb3xT69nI
mxY3hohfvk3okA2M7QDT5Gpisv5A8CzFqayccEgA+lnFzvbQFeoZKmAhAXwz+f/0kkyq5FlVZu3z
Zg83d0Uigu55GRC7tf1FuKqRcfx+d40KlRgRoAiqmyD4DJhoV2oFD9bGb8GJzWxFlNWMNm8I1IL7
wSqUrFSQiFngofDvG7kVfrOyTKWEBQGvMMxzkc8gzSRiGJcV7+GIoawKhDL+YY+rdRNUiuJxZRnN
N68KeOtO8k2PZMAqoCIjlkjdbBktSArhseWU5/yB8hjnZoq0HjgRjAmiLRegVSPBYh5Ihi7EfgxU
uuln0Ca9sQdOA781uaiGFhShrOySymWidoOgPnnRlNkZ5MN2VZJerGIN7mt9FIwrnKxh+idTMPxm
rzHky9n0ZjalNtByQM3o+7nQkrv43TK31pbJUaMTLdXzDq2TnZ+yzyOFlhD1rfZUXRT0gRgFYXj0
FWAEX5DCXAv2oFmt6jPMAqvpx6P1wm9RWcI1GtMFPvt5xZ1CGg89Z+diITa49f4FyVeAaANBwnXH
D2EPmMZuT3Qi9S83T6kHtzDmLyVBAVhRPvVjrjvHw5jcXQBIIs4QBHYwWaHMn4Tq3iXZx2i9uGKn
JmLtOzvxr8E2zxCmh1SSILqEvsMtnJt6Wfjf24w+0brhi1q1IRPUJ/ilMfSqhkcVG5m8qGz2EntA
l/9h/5zmsNyvojwMaN1JDN6S0f8ZMfPzMMax5E0Cu96nm3aqq7fsIUpzEwubqEnk7huya+LdH7K9
J7llHyIJm1XRsYfypedivKnXSCRleQLLO+QggNtwbCwkGAtR1SjqvqnsXYA6tozP3adco1cgHUCF
5vBgc8wEb9Y439opZgmnID7DSUWnf/UfAwh9KClZBHi8/f3/fxZ/w2PJNsNZufcHLeWw1Ic4rrKY
lfbw//ZdImZUDcxQjzUZpon8EvWpD+uX82vjK8gPZGnIQ1yLCbVnyTgiVGGZXJ1L273daJ9Jo4h6
Mqgu1a5gzUSfLkz5hgZtUoLha8c6L12twAZZphdYNAGD8Nj95X+ybV7yaHiLtQMvFqeaVomFrtft
mjoeBowL00RvN4rohlnyXinKxNEnhl72xcpzQFNqkkckjzt/9qOv/98/JhxRwPAIfJohi+RTwkBT
HzOLu3iZbvfkcgVFcEwqPZnVHcHJQmMPeseya6Nu2udAF9hyG22hwkbnBQzvMk6DHnrD3jxOpuw6
WMRcyCRE9BkdAyBEtvUmP1bjdNgFFV/zPuAF6+SfA2pP3Qw8pWLGuS6A44arLypguoe9Jfm8ii9U
VUrcRvIEbzNTrAoN7PWM2krDAStwTe2oQqJLuaEywhajwrIXeQv6Pf6TSulm44N4m9vinHEALupF
s6wuR2m4t73eOZzyXHxdH1Myb72S57zsc2cjqADrTUCyESR/W0B2DexIJSkNGt6lMSDbTbC4+1A3
MzGXfS3BaV9wzEUjE23JbUNuoNX9Xx2smt4r3q0c5yY/7isqA3tqzMsg7uSmYoJF4gHbtsquTmEh
IEqqdGMHD7HfhxM1n75R7eB26MqGijQ5A42GuVVLU98BCGK2HaQ0RrClfqCZFnai12NsU55IU03R
VqzPUGO/0gtYV0HWCya3BFUN/e5t9Xc2FL6UMqb3gXXhNKfeKUh0wNVwAtOp53rH2gKrm/IBNedt
iAKD8c8KDQbt+lpAC9XwvqpOFn0IWAELs+EPsPl1NOCSw1dmMtTRKYk6Y6atCpR7w+vsWW9R8Z8t
fnZUYdujdMfqeaM/A4gYS8XgdEyKpB+XnBe4BQz/hnUtjj2pNbgHaPx0sXAUCrlr4CHytVK2DS8T
MhIfwT6fsLsohHCmOWFX/Nfh8X8geZPM58N+RrEKaQ3Z0eJGGEWwmXD7rKN/IyimXigTTqWq4CDk
UNpviWlm7U0L+M3nCFwoSMwkdj9DB2pA83gPrNNBPJMKu7GemxpgoitPAEX2EiSNLx/K6RVZUUix
SpXj77emXK+4HOSCzQu4ulBeqQFmdpn8O5qNZqONpN0fsSRNf14iCg1MttYE/jeKVhqDVpyZiZXI
3NcIC6Z/dpxNKdDWkEwuaIqLEUpnIZ3zkzXO04Nsnlv/JmlC/pEvquXOA25KXk89kzhdY3/K+C51
O6aLHKKCBMBOk8c4UWgVIzDF6ZfnLguznOPqLOuh7WL9oJd0pcw8plFVW5C3mzCat/5BNza7XugM
uA9fvXwfWwuyID5gZw3bYgbSiRWsdBPDnjMA6UurZztr3tG70EAeQUceIPwGzfvewdmb6BvcwenB
tCGpBZGfzo1xLGYxtWhHmtCAIAY62eLK2p6pTJhnDCSoKezFajdoj+vIoTcxuOZOiwWZpADnQy7v
+ZOBvq0viC0MjZNGQH8lw6BVnB3WLG/HKfHhK7lTYxRY5XUPpbLeuKW3waUGEiNsJ0BIsdEfR8rH
481wpKdLOJ6O242NJgeUkXKu0T7Af850LKfOn8wYn1BW6sY2o4GYUjnL1JrYIp7A+B5LirC598iq
LA0Yi0VYBDTlKitcUioOcM5TrPmgM4YVk+HMNgQ6mvkGXVSrIBUoIkmfLH4Zso83ItPSlmo5Kdpy
wAdKqU9wjX/7JdCzjMus4FT2dJJV9uoTq6pNQV9w1TMdPvLUjEdrQmHywmIeuXjSlwOSKjzXoTXn
t/CCRegX6ThHmGNfTdSJIukPeBs+z/FxfCHLTuSqMOdl8AUIqveZ4NwvwAGMHKIqkEY7oYcnLQiO
5hoB1bjNDePJOo8I1Ltjnq8qdPnyeYr7QbSv0gP4SNDUtS+DRDVG3kVfFBOes66xO/iNRPK53YGR
gpbD4x6nZ7PdishnKqSYgwhEv2tEhXbJjr1vJQzqoo/EVMhe/tolj0+Jw+soRpie2C4I/acx4zb1
zx+CXwzowCBRerTiX55IVdzLdclRRSk7k90yWvtqG9VaFAfPC8SXP53Bc509tcplmzthvwZDoPjs
7gZDhwfoLTRyvTORe1+J/w6oaCnD+DnIC5Xg5Bshlmq+50x2riIObemZRP/v5WmbfbA2cGCg9IVs
ojnT3M5YsRT/sEeViWWcFv4mI7/+eBjMhUWL5V5MfqhvSbAfwTM3g8DBQJmPwO6y0sGmbYI3QIK/
KIOE9Td3cV5XUeYlYScZJFx46UiJS8naFr6yJwQlA4Ze2ltbnB70S0SHuKeO3j7sjyklBk6N5Ch8
peUmJbVBP8m9uizX5C+Kjl3nyNaVzGPtqRhyOPSuP22DScp/3vY2WgUrJ7lBAkUPoCzKantpvfNT
wIjp0YHGkwAkRG9bj/PrAkbsgFXwG0DqmHrwImBQlrB2IFXkW6LWn/J98klJVqK7YyveXPKO8fBs
iX49b64Nq1RXu0W52jqVBemlXNDjIlBA7hQDRGOi4zxIjP6ioWfY360BUCS/hYfmARAV/jtiuVWp
ZR/opLLmkL6Yug33w7wsHWh7QU5E7EgA1XtfnT+oXeNv6wuBB+XNpgQ/iu5mTZRmk2Bl6TlwJoxx
riov0He+FJbiJM+4Z0X7t6YXuvUAkCgV/Ao0EVWp3JvzWOFiDiWnVGbmELK0DgNuETAB9aU96Ow/
+KXBHNwDHj0vc5/Yd4Ad/94yw1WNcfihCOmqa/4ADq0I/jHYo5yUO+yRgIWf4kL0HmuKD5NClwfW
9g2U7OTSRJaYI1QgGTSej1Z8gOXccyFA6Rt8Y++8mT25ZH3kuEDj/nua5P5aiMq7xe8YzCgFn9ex
LQx7MPA8gyNjsnkj8Mr7dxIHghP01NtlYp5nC8aJtCn7IwSIWavFRFfCmHxpHS0xFfFf+IvnoGtF
M0kuijiah5OR4yIuOEbsuyz+Nnh6om+NVwvdAVLsER5FP7r+oUpGrHFYiWT0qq+rKYlZ7xXKDcLI
Y0TeUuV9+QBKxj8iV2c48PbJgCDfMIqOV+9L58AmBWC5n1Fu4n5GKj2sli5bAsSk31wAw1YwZAMb
937tLi7p1EEXQmMCl2xihYxx11LwSE1LuoTCxDQRWR2Y6q8n8tXKmiE8f2JYKiercA/NDmPu1HZ0
2XIrZx3/JbLymgf0u+8C0yxnVQSAAq4kogqwtza8d998X7pMiGCYXORtvYaW9Am6YS9NZmLmhw2C
IEjyirC0xgf89HTth0EygqPMEGp9S8rmBNjpCU5ZNbUwFYbBJHZ+1yk/pA5L00I1NwbZZkCIEZUG
9FOLre5dwlDU8c5W82lGx7hs9lql7XYHiRsvOkeqVmCbJBGvugpeovGkwESJRPykShmpeEQCXDpx
U5prFI/y1XMDnR/Q8FEJDh9SuK7jbs8J4qK9xaC/ojZEVXir4rwWfn+cOWC+2+LsTBLxSEOORkoR
Zw8HcEL51NRZNv5qaYNSvaF4bvbVjKlEPKxToo2T2y3eVbd7WGPYoeaHEfo3/lzNt2inJRAnXt/Q
Mdu9BpRed0WDpt9y+V6kYOJKgA5sSfvvjKVs6Ghc5AENckXRKMxNqOOTeFL+0yvVjbdhbZk842Dl
sv47vMHCIEJ94cvwSszVqn8UmpPL+GLSoqauN+mTNJ2A360jALTZcT2fW/lClCd3Z4RN6vLPJ4su
MDckppgTnfLTokJdmZScMlBf1yspxHYaFEk5RnG660xx+RpV8/H7qqA9fZ/2Uz8G6r3Jh/BAF8p+
yITzoYyqAo2SLKEcZ9Pn8+7NQYCw9zAD7revx+pWkzRb8hj32YLVl2a2bZyjUrCcnPOUbysD5ZzR
iJWmSTJkqFwd3dWNEVw4czS5z1r67apNHXCEA+20gzAp+5ZrJQUTxwast7DLjavBtTOaSQ2YuJP7
0eHS/p5q7EMVBvCI43+Wf8P2GdOQlgE0x8vvZRu3nXBBb5Bu/5uF4w7126/HfIVnPthBphEs+zVK
LLwyd8NZ48pB1BO8TtZ1Gjj4mthpgpC3sk+F9ncMsJeR7rQBQ2VRw1czDemQg/doOLONQklQCKR1
JSbZAkwN3OK2Ae+wr42BhH3/Q/6B4BLqF+Ulmy9o2XGitjiw255B9Y+4xjhTvyc4gfb+WTlhldWs
3NDztUuecay061pi/pnwUlbba+OheeqONgU10/ZdF4W9zUQucDwnwBRnR0Mkl9IdfBNTybgwbscA
/3A3DErNSMP0I9atdYAuDUUZCJcLrxY0EUdAQ9PF0QNMGCXKbjzTmv3VF59x/to/bNfFZFx6tW56
qB6lE9F0nBcxUeJAytFpsnvpwNBxCYLYgfm31hOj5f9EvTAgQ/3hIIEniAWvOW2GnhZTDwPc2ZhB
cvTx3Uovv/sdYe50beNKPNA79NWBPU31mDl6endaQZ0ZZ6u961FQQUfXm7xQ87Pp3NfgvG04tXO3
vY4fMAMwy6/3PQJG6EU3I+keyvS3J2O9sOBEu1qJCPmueHu/jRJtKavpw0c2SLmFHHmFkxC4RRaN
XY0VKVnxZ15CHDlykCYIj1XdHGNJaUGrvIQ/XnZlv5cZTI97Ln5lVVAudWtBJC9pA7EIPJOX+vI6
WtoRkjhaGQzak1rLnQCMUFCj/7pfLLWLMwMjBPm8a3/Z5NxvAG6mbJVAVKrh+oK4KBrfAZNWAiSK
x34kxfz1r8rjm6yR/s5l8Gsz+T87VnS5q92B0ZOjejAcziMPaN+zT9Gfpljc3HWBAvoxU5T7JSka
qLi77add9JB+9ckUo8uNTrHp1F0gdTjPQD2IUy3FQiutBZ9nQ8TMTZlxRRT5g2nSHxWFsjEi8Lgi
O9JSkZP/QQGdw9E3XjQ5t1KZPiWuTfRC4m4KT8yhgkFgMr1R3Wfb8TMyVEhRnZWlYPznXj0VRReu
XMKJUTyCpXxTYN9RewcKy2js3WXNOFgXOTJSMbizMApVig2SacqlIUNWz0bnDX0GYPa0TZH4u86l
a1rgmORq0ux7cURH8S2cqGSlYCajLui7PipbgXC7cwLBh+B16ON21uQKXPZXrRJ6I7fs/Y9TMFRP
/YiaYxQMPX5weiMKJEISnPTFzBGzQilVSbqyDsd+QgOSbkj7fiGSP5kCjOcenksUcDiwy+0skNor
sUGwHQ1L2jdF20o0Iad+samVKnboPQWlmxPXTaCy6LlSOguMXwqsyp3CNA10FFzNxcmmbwvBcAWS
vtZ11nWNnqyc4UK+bCZCQI+wgrBI4blYrM7M8BzGnZRpQdZhkfIUq+YKTC+xRkILqA0n8iSFoIVG
vf1dF7rn2WylJzVpzVSJtIDAPSOWDYhJ8VOrh8UlS7XHh53zjtyImUWm5IpbPBMlfUM8ppGsrmHY
I5dutg3S3RSxek+CMnK4IkSbyX28xgTLmRMenNbEUcfvulcdI92aNAtCYMmVeJaqQko9v5SuIj4R
x+KeiLs+V7YMSSZMAhQ/wbHFzi+XTNCqC0kyfgUbNRTeHqeeveJrpesSdgV9EofRrA2duRmD5uBi
xVQ6vSrYzhIuevoDvgNJabiLyz2xd6Z/jE9R/tQ9WNTdMjViLEiYylVpS94Zu1sZ+TV/d/tqv/XB
vHBDBCCQdid1EiVU84VAWSZqxaXbz2YJcqcNL26nepntl+wlgBcaMpLdRJw/85zvXP953Wf54IoJ
JsUqTZy1yJdxdwUl3AK/gTYpPZLRa+SYwe6koYpkG+QflKVWYXojMkNdV/kb5GXcon2qjOpvVaSl
fXHnVKxEV7AnpRBVDk73N9fJYVpi2b1lXvQ1kGRcA0NIUMUFt1U/7wB/Mv1LJ1bnMDvWEDcLHToF
C5qF64Zxbiv62qdQNuwsU5TlVZeM7bkGv9chz5lIq+/CcI0hihKWmvAiCLBF1p0hAeEh4PpOu71p
Fa4X4FmDOO1j2tIl4tNQNDcVpkFwpHeKbIMdCVNOf3E3srrnAUqK+lL0b0HNe+U/gnebEvJbNBqG
LE72FIYOM0Mc9rQKCudV4dHzCAYsrbvG0GvEcr5cK6C8haxUJBX2s7RIqn9iAA9jGhN/iKv7fCoM
RPtbFjrJlcBaVEX7q7Da6NFS6S1zoOp8KPEqODdAXHDbdhjWl40JmLyo/+G7/OvMuLQ306dujhxp
l+pjDao1IZuCC1s+Si7uAWZnna47ca+Z1Oog5ClFBGrlqcmpPhBi2ouQV4nRQzA2/G6lsAJGixUp
l29f6OAOv9BGzFdI3xWWd40Mlr4QSqipx/EaykeOntaiBm1EjvcTZ4mcxVLygod5jXWfwuyrWAjb
n1q8hQUkqgIQM92RunydCQIhnc8KzokuTeGDSAq9NEIdJq+8MIAYwyO7ZBL5kL66VVlSS2kSbrYl
DM51zbji5RZLjfkil4bRJrDoQvsdSLm4JdPMQmV/KqnSrl334xbJu0+6I1e5TkqSKTN4jVfWKZQh
VrdDG5ACI0eaq4S4SXHuYC5vQ8ULCyccPhE0KnwskShqrjXoHDu15S0n2J0oY4qmxQ87wnOfOC12
pRMYortq56cc7WXdtGSbXt1xknz/67FYas4UQeGRRKEdl2nfkyqn5vCkxYImQNZjhyJxndyKnirm
GifnbMHTCO5lStG5RonHqqBrDX2ht5iQbJDyGThillEQCbpDiqVCUTEzsTdsIuPmZept1ch+cZ8r
nDu2xkukViC1WY93C4VkAkxxV1ZsiNL2o/YK7gVEoD92Z5+h2HE0AvplrlnONA8zj/n8T13FGjj/
hcoUObabFu+9fSOanAPSzZZrcHXPEULZtLGI4u8qrtHwpjtgnCnxPcgfghQb8dJjPXIyorSR+LES
w6xu7JR6St9s+ISI9FPCODzcU5/ks03p2HQCx+usRS7kZkQojWsEJNVH8z3z3CQtvPOFpthhg145
0/Owcwp4omhsSouK+Z1WwTNBlUzwtADIsMlsflDZQXZMANJeYgoZCjwG+ZSuCO0qL4PfINUNhz1z
dNEPeOxMriaVu+mXIv/p1B2UCtnyFr9rj6zob9Fw/k4LhBcjYXn1bES2boG16x4fXs/VcflbUL2P
Rm+reZMPG+ELQ+oGbAF5LUeDMnU6v3EPw1xV6zTMzkEC+/qJ+JWRPiIXPZ4jSGAlXOtjzyDuj8fU
8IFplxhk8V6p60oKE12lpZH/rwx4vOrsGybp8cP0tmbMkDOhBRHjlj56Yb6PJXhdJSKYhh68Fjsw
yje7cYVY1xRx+55Sezb8PK+7ZiA7jBaanlysgDJsQiEHogoFSSowb8k1n3mGsuC/w4i8MSAwdO82
SW+nNXFad/KqtpA18eoKIiSKZ8gIe2MxndAYFeyc39PN1OH728cvEzlm+cbLy/moURftCJgNQD+h
EX1BT4vJ7TtMuYlXMNkNfrVfOyzqpmPlj9G8r3KvD3SwUJ2UJEcvb8+CReBCYwmkCvwrGnNx3zbW
VzQOkwthf1Oz4M6Wz7BZ/AdhWUHvYgFovVKXCQ3zX4fAJROH2lfp4ZbiF23cfxJ75UgR0DQdgFkl
VAM3VZyRB9CVgdZwPwqKtZuvrWn+JAzpjRdhSK6HoovLrzla79OmnrHIf8/y0X3w8HA3etPbzBSP
axP9wTUddm07wBrwwa91sQxR02Efmp1z3VSCkYSkTEiwQ5kMbm1KH0QrAlW4Z/I0CR6Fogq3KGRz
/Xd0mRs5pFtx6PVlo0JOHRQs6bqmxhJtPMzolrpy1oCbi1qeMuRqT45yc7kiv4rlXdFEzaT1UC2z
C1Di3eXyV2SBFpbtI5Rfej8YizyjWrVnOeVj6srmvf/zxf96eBKUG26qmz+36BmFHbE/b76Lsk/f
icdaUmqX657p/mNL3vwYsxbRP7NIeCAfuSUPiKa7vuxRSaOUOq0Ljti12DEM4xAZiNYE37kxFBx+
/rrClMpdUEwjLPr7xSn84ZkXWKwcDoIroNX7U4H2YGZJpU1tMYHfPN3BCXZxp0iZ7SEOnV5yGkYK
vghDq0PqLb68JE0CzjegD+NxOdStmO+ElXu4UMYMMAunIwadxiW6YL2Jm676mF7Bim4ZGbtkTRkI
8v0Y9nDuYSwSqgDuQx/76YIn6E4ql8cxHjAzSyF83HLl7SC58ogv/e8e6eoA/AQUW62Ce5eXHHv4
EdykpiaQOlLwRp4bkKXMpKlSXSaDuVNf1VRYwxQEcTZpGRDzxj39b5Y/RY5klaWkE+l1k2KCvxLl
7DQRZnE43x29z9Vcqsv9xfWVTyZg/zMxhaGYhFS9EtrTaI/QwuNXiUV6emnboLPyK7Yc5K7FRtKa
Lmrb5AuX0EXfyhKA/DaHip6e68xV+Hp10crQwDwDLoOVAR4HLBKLMcJ9zUPMdWoeG/k3Yj4t5z4o
hoyZtWdW6o7TAnFYT/gCLr3PaVnTHrCA2wYjDpxGxWOmxuJTHTU7QiyqrwVizCID7eHNKl7mnwaV
KFdtGxV9T607N6B72UGivoCPj4EnSSRBafiDKkPgsd2MBTN+K+hkxOInJCRzHPqw7f/N3UkRKLvh
84/0jcD5ITDtg8l8t7gFEYCwf4lMNvSxC1xz0q42qWxHRFrPMb5BhYLvmHfB2olVj/FnGGz620ol
brXEyjeyqJ9mzJb0xxmObAlq3cq/JYokcJOeCHkjUPSG5BuozM94nMFgN5IM8IoDVjTGPKyf2d70
XPSPxcvwUL+Yi+ERmQrERg+mqXR+vz8glAnyOR9eaVr4olFtC6zUz7qe1w81FNz74jv4J8gY+SnA
GxuaxG/u97z20X3WS317JFcoHOoHBn41Fg65nH7nfAyltPyA/xX5l6GAwT8S0vuUdZpZsvuZDEAD
YQ3quQMQK46fAgopg7CPtYhZmGlv2Wi5oDSfLMEC3TQnzA4Q/tZxqTOTMq/4/c3GdWPM73OBXNLF
CQEBCHQGB4Nw92IRtHnPejdejYVHHVqQJLPKjxJs+bY0Eyq0/ezQC7RupAVwKK77onuMT48phyh5
4+559kgM/Rqr/NV/9cY5q8bS3F8i9mgwkVCWNmxxlIRSeyWwHOmWKiP0yeSWQOziHlgTmH9U8nXj
84J28cFDIruLmwbk9BDgrwjXrfvXAHUPJo3eybB2OQbLQTdmWxwvdiRiddr/Vxy4t3dYBIQxerNS
gSpjSofmGHXTFpUX4raTnk20LL753LJcmDKWdpqOZZh954LK7fyFkCnR4guOItsCpW5t2EbrUqtx
rHAVpLbXRIc2xT4ljKlRMSYHow/fmSsn6M1/7qmdZAx3nIoLP51bUP18P6bCMM21/ytmYhubx9FJ
fZTbNnZPj5NL9xEjfm6/EKBPv3f2ODNrRTqQ7+9oznOH4bx6uVfgw9GuW7LDed1V+xW6lOvnUKYH
G/O47qJoFbFkAqc5z8TFmsCX4MEhgTSRwSajt58PUrc7JnH0D5ddcF4re2pjo+COQE4zMuqOoT90
jVfnqzOnu/96r3SWsuA2HZMHjUKf6seV2ppoZGMGxEGUAwTDkXU4eyxqKNDFKi3sFhhGAomTF/IH
qhRB8MDDMXjRF3mOgN1T++xN0rbMW4D5G2tol7FsGuhnBenv8I7xkbdksxFrgt3skMK6jcaCHe6W
UK7Y96egnTCWRyGQw8gyDvXXK07ZxYyd9aFxwlMHl5q084rTKj/RSgNz3hMnyHckrSjuhiT+0lbv
CcBw/KzaOQ4u/ccwrEwrVmEqfg/cW6b+NWS6xHdfEbtP1UNJ728z/INWddndO306hMF68QRtudbf
qei6D3fJtGBSQz3ejhf6//oIJ32ua2wqRFYWN998W6l+6/lRTSIBrBJEG7RzcnUd2YIj+jr9RSKm
NUvpjLLQSVMdtXZ1JFpdXyr23SNDqkhKSwEmZFTw4mvJ4LWnCIYGh4vrX9hIoaV/W4Bm1HThPPmc
m3i4XSY6yJs0Dt8DubDuptvZLgN5uh8B8JyyWLbD/LNUTYARcdInaSt4WuGPTV+SFUiAA7EQdOnx
RIpbPT3OrooPyVdsc9f3ewRSLu6nOIw9NZYBldd8Tp9E36UJKAbmIW4/ET2l0AK3e6yG+MvxNWCN
+YglNDCPUmMFDRfaR+qGQKXChMsko/gQofWXyyEB2gqnMa21ZEugi0KuSUyMmG4osAS921zVB0gf
GzFB676ugmfa3EHiTr7OrZMozsQYdCdEC8EXaCzbkNYZKOc9uxDIZttQ4rQiWwrJZdPovScrymgM
kXAf7IcjiRlPY5mQ4JKSej1dA7sDw8BXx8xeNj4xetEABbZprWXXC3Fzd8fM0LSoCY6U4xsGvTGq
Q6vOTx91L16ffvMgLChmGUMPiBByleM6ZCBJy3T9aC68IZ2ghWi/gJ6MbPhERsVB3l8lFnpaFzog
wZnQ10hgWT5ovf1k/2DNbJLFQVWKe19fsdgt7Ji4/hzbM+n1+fwnWfqtWGebNfowQDq4L3S0uI5r
X4cl4ASexZinGIeW+dfbxScArUadC8QAFP2dukyqMQILsrdZcMZ44YIMvJTw3E+XdJLIg0xU/UPQ
MIa+Q2tk6FvdLILO3zjxgAEcS1fIELr+8meiez7NKlfzKnK6OCjxel6Vsq3q/yqcbrAaqvsQOxOE
X2iISO6pyknulYttQCNkA5gEHX5iR/j3X82ehvs3qEOy6hcP2ARl0EvrrdHYh5T7kbetHgoZGCOv
VUh1RucuvOPPm7cpkTvdeYpqACipwQnPC7aDpNMKblpAF0AtedC4bFJNLVoD08aaQgWdEDMVIi+o
oX5JyRKgaXwVIOCQC5CLiPMeqVjP8Jw9k5UKH0A1FuGdB5AsTTe/IVbioBi4nnQirvXIs6AHMON6
SzAMTwhFvEzxLE7Ev5Do39Garl9V/gNtJOsySNvKaVp2Wf0RkyFF5Ivyir9lYL9ikeOeSr1FWGe4
MBaCRwAuetDDvtJ90ccgCbf6OFNs5gI1m9yFcMGvKNXZAj2+Qz5EGXNDkwknFhhdkHqUiKX95kY/
+Ufbf2w0Wyw8Tb+HlwES302xiKb3F/YcWIkj+942QDXWq/JGw98pPs8bBQVNEbQOpI4riKJTLAnI
nmhBWYGsAY8jE1LkfjUn17U9IrmbWCm4qbfTppi67w89HaulqQgBs8/uqUJksD8u+shIV+TLbNGx
hDN2rNK5V7WwbHHpcntUDSArtPz7mEebRAdWLrev/AwTgXGhlS7p7HWxW7iggaBOY9FAbXHe+93v
YtMJ2FDu2gn5JxU/10tF+3vn3Rdh7D0PIj2DLt2dFOU9DYYXa3ZkYoxU2+DHw/QtLtVz+jLKVtl0
6274MC3fR1CCWnuRFDyF7RXAELGCt5c5XfZHjptXq29TC9iigeHhnyNeVsqGBWws23JuTvOqc0ud
cw+CHnCQCxWRb+93Kj5VC1fHR7yKe3ej1RDwTwoiS5+RFt0TMbqAXEum4YRMnEMBJKFMlAC7Wmnt
Hjbg133oikOhs+qRPo2Kh6vSlvmkWoTTPkewmio97zZrHsF6MsBML7Ov9oWRCdfju6sPL2CiMzTQ
XkgXEwLxZcYIrHaZ7zOTxTVcxRSCj67gI81V1bZPJSvz4C/M7D2dC7ZF9F2q0XT+MhruD40nX1iI
rnJABbFlzR5SMEffgdNBfurCLMIwceS/7wfWVP7Ba6g006eHk2UIjNWRA9ZB0RgwJ2F+L21504th
imKU30wSoZLUs5ApyZpjXzyffGJxAGu0YbUHVovgUMSHC3FeAj6E2p1HpzRuX84584BLrO7sPMVb
kwFodJzokd54neDag/XWzYL2a8I48quECymyoorfjWkyk9FDvwSsJEF5CiEu0M9oLKaREWnQDZg6
LfuTrQikh8IPBIv+TMdYyrSJcmgwLVVRgNF130gqjd5tXL2MTuIhMODTPjnLwc4Q8za2lpwkkRk7
PgzKLUKvE0sc2ia/anamztgEtXeJSNkyzdXbMTMODQNL7VS33m6AtiuZAJJBMbQMzY3fpbxP4RAM
2HMpTEL76kIhz3tLr8PdlKfaWDcAWD6XxQwiuuadH+5YUIKxVd97ebTkiNnCC02ipqkU9QoEGOX4
jtu/S69Pm37dQ/asCH1G/1st6Ka/pDEFSOg1SKVd95Xsgg5I7gCuaqosxx367vdfV55LL6bsgmmA
uLTdVijp2O6aaYhjLr1TKxFwFUqfqq3CY0ypP0c9PI8Ojx66RWAkU8NQf4UHCkDgJFqWc7BlENQs
x8IFGll0QO3mI+RmiHTxgy3gzVJgVwC0QC2j4p+soHoT6RWlXuKZw1OvkqD+/HV2xVsquzbu7Mpj
IZYJ2SPYYuDuceAovyErq6KX2T5yafSUgO31qR+7UkRDXyR3YJ1i0DdbslbSv9pnCnN5lDg5yhaW
KeYMkRpPdf/OiQEjODCQG8kvrAgtUBZ7a6IjvpOLKgbmDVvw+2ofefM+IqJbWrr4QVE6Yp4F3QLM
cv8ApaUqwb0xTjPtGGcNDHTm5lnBs9W3l0DoorpPquizvqCvNlxlSqhNMgk+LC6seWrwMOXcPgXe
a5N/bKPUjg5LxakvSjGVMShV7Lv0kUYOToiaMY4g0ruy0rxpvpVAZ5SDCu8+YjSxTGE1dX8Ym7Pm
y+YnYDx8cymyAerXhRFqNi6qdAvlVjIbzqqqkxX6SevYrQM8w473Z904X6jwLcZ64DCZUK6kMfiO
oMzvYB8NF26BsOanXv+opUjrjm1MGh3TcIruC3Bed3Rri1lJFPjKM1oS45lKSP0MmSo7cshigE/h
1xXqgScjQtX+Aw3IOV2SCOsR+L1wuEzc1Ne3iRBXdxXRBnezPXWkx8xLz2fIAZT8fv8AzYQxbCBs
bYjrRhYmZ0cmD3DVwxuP7MwXewM24VjXtxGrr4jitNu7ONi6CeAG731lZ/TDwOxGwaCi1WpxthHu
06SWgaoHsRNc3/Ar5yy5UUr9RosV9Bne3rXfiSajltkANBhMSOVjP0NoEaL5brx9mt83qs3Gx7B5
oeKuRNAFJ4QWZiaHn5eKHSW1f0runYNSfQto3qU52PC6z3JZMP+QBx6+hrfFNaDjnkJxB53ZD8Wd
lkxsSmMt7mQe+NMW8vGMZGGsNOpeoNIxconsLqF5nlG1OJSNUSecp+H083FvUFLQtBuHVbk4wtAE
KOTfRNSWFattYNrIVrroTyfmiKheWsBj4V0JjsZ5Jt5OXu+T+b9DiqNoP+cz0caQZKVzSQ2N63WA
5JDqXoMy/WHtUiI3p+/vzFXLpBWI/khYxxzdzJw2gaiqHhbLZJ59S5VgLYZ7QBghkVWLs4BNNKQy
kglIT25UHGQOI91k2ygWtayM3xSu85scyJhchfnf7QYwLM4hxo8TFNCrgCoxPYF8pwPCODnvDldk
iVbIudlQ/54aYqsNOxkYAHHYAQw1k5MGLYAm+J88dAD9pvYCDIESeXdBvY0FPrz648sqn7gt0rxO
z7diqfsHhNyN3F6YzLCD1YRgjRL0orp/LpjT2/9lsOdRoxuGyQI+E1EHHvSdpN6BAFIGVe1Ir2Cj
WzL/wdCyglM8/RsxNCXTyFVvEq8113Qf7I+bk+HWbzhrr6riogOvdT3wnKdJGdZfM4hFIsWP/dvH
n1IvaeKG/otAxkFoyoG/R6WZA+qDtUt5fkz+biwZxMnvKnnbnqVRw2V7N5/wBGZVLaOpyftgNzGm
k+IZcV7R98Ul+RgSPzX45+pfeTLQJD46znpUDV4ck2B63wBvFCwOHf+Qu/tvce+e3y/ccHOVmilC
gR2E0HfN2NvTakeqK1QyBoS2E/H3XRsDjO0igMrcKfb6lMWgDqQaDMarbzeFLlyH0ADhUQO+pyQw
kglHayMCIOGGW33Ug+PLuiND1C2lsc5DFGPToauVhg3WAVc6HcjD8CgnZ75M45JkMbofjTLxTwN7
oosOcOVOUWzghM3e8SaVJIJD2EumetoL/3B4LW4CqLhuowC9SJvGy1rlCqvs0zaWZ0aAm9fLQJ8N
3l/8bLZ2G8cbRxHohK6/NLdT7mqyzGo3smRF3FOFJkLYCJjKS7PiUkUeGjFD0fw5Y2EuU+Y+PIDT
qy+rilmtpslvPzoEo0z/eiFw6YpkW1AHYct1YzaUVfUiHzewktiXfNBttMCG58lsOWQRpN/3y7Ic
EJwRkG9Gkh49H5bPC/pl+DYmFP5MLawIHAhvcBioIiTv67S/0e2Zc6NrkX1+Ss7DZ4sX649LxylX
vJXEzfNk6CKJEq+fLQxav/Lj8jR2lgaXTMb8Y5vpfywn/+KgsRIXLaCcMHYOOr8jMUqfEdpwIDd8
c0Ef1YnU30el0WkYXDYSHKmHJCa5wQ4BSy1nT5S3JoFsM9a8OF9NGUruFY1T6ukEptdZnp3m1rsI
7R1FTXo788/GfiB1ivPcl63TcCAMKImbrDp1E1K1E/jQi0VPcb9NXUxCEN4bDkazsxPkfu5UifPi
ielDenvxCxVl1F2nH9Ze6TXzMZdUh4dtIZ5fPECeygWPjXMU7Xp9KNjccPJSycDUuhFckHaJv2dT
P1zaNerSv385SsUio8dcfuZfmRsw9EoKYtjeqrLcXySiLMgN9EoCZw4oTxZFP7OQGR+pXA5QBfIR
U6iMLinrupKYIvKWlIYbWPn1yNq8j+npvLaHsjOqyRl/G6hDulKdNLFTAB6YMDhU8p1VidJqeEA4
GhszKCpGDG8aNVjQn3FeYDhgrTCTwADlre5xvNZHuSP4RpUitIHYat0QT8y+XM0lfwOLSpXCduzr
GVa9OjvIhxYKvLNuFJ3G+mwv1dNRPKfT4D7Z/6SGnqlOKQEgkw1W2znTLBMcw2qSKQAJkNFKd/5g
Kd5LUSiAHBP3Av3exHf3IMpZtsYspBeEq7gU8dp0OIfsRfFNnMlhzxKIzxTlSosCYzk7OA0vGD8h
bijH2UYakdQHyuKOhRbiWmftQsaAdlpWcM/xIU4NPrTc67NoKkf7nRPZYxINlNbYNu4wJw8lF843
qfSj1XUTh0fLQWmDeTJOGcUqhVPaL6Xu1D7snQzKElehQoUkuXO5jqy6ht84aiylA1N3Ysd9+nup
aUv7KNXTO9jKAr7kFuIBt+qKL8/QblDJ/DBd6Cp2OfaudLclg5+zrHgFzGozBwN3v7mnG3UhMCmU
CimWut4kNh07Ha9h5tawHhoHOrqcasG7AO66a7HgzSUalXeArdyMCLPOzuXy2fDW1obH7y5fShWD
xegSqHNBabhNkiS8YA/rNTvWz/RCs2a0WCMYbk6pwtCOXHrfWLi2F8OFXQr53WJ+zz4OjWfd/Bcg
cnZO247jgBCZwpgNdkd/x0qUTjrlEZqFLRT22pI0Jy7MDFvjrRdXgnRG0zQnNnzER095UY6dgvlU
0YodjPTCDqabm8f4ry57zN6tbT/sX0ONA6+3bVAScdSgGfi0r7zJLbemXgng0RjMhaWSjJI29QgN
G1TmdzuJggwF2dTSSCbE1oWBpgnjQYAw2FBswHtzNA0iuI3jZ/VaNMx8CpjcF5QAiLHDDX/Plh8z
3670NiMgHEIzpxpdJQqoV9pYIel4VD4hrN4Uer7mPvYgt3ZCYaUfz7ARgcStusKvizqZKRxtsHca
tF0DzKRJsUvAdRv1kadPrYl/HYkVREGKCeIwiYaQdatzh+yj/3S9oGbIIFyx2jgZ4iu3jjr4UwUy
dLbFXQ9sM/SuviBV8s7hP5InindFXaiCPngYzXUm5JJUDcx21Se4j843W485nZFMiBUv2dr9tbnC
g9HkONrbbNAbEZvI0V2jTPDsBn8+cKmWl0RS303eYVkyZhdnj5bSLCytZ/2tiHnynwb2Nw47Cm3N
0dVIFNSwW3TOrO0N50VULQSdT6IwEr4xLCAnACasSK4skxGkGiTJ5w3HUfnLEOLOHIsnc8H+/zvR
MAhhce9deQ/0yrT6nsh47tB8fY3q2dsjREnffLGeM2z1s0fH2F7Dho1Xz65ozSySxZ28oPqpWuEj
oaLfi9TmlxMsiAjdWlOM/GU8pog571ZbLje/qkYwa0Y+xjYzhPHRXbWHK+TYwQrh+QUtbr1hRNmr
hn8i8NWYH9lP2eT6cr5Y3GsmbeKj0dFphvQc9zKkq/O5qTk1XQzymt3ZSM+dVcTEx9Apwd5DxzCA
j1v9fIIF6an/yoEynoOIdUPYXuwCrskfPka3gqF75VaUmZT29Jom5QQbrhm1cOJaFN7QimE6/l30
H9wxUErudb3aC3O4jZuvxaVyX9Zzie1lwoWZ4HrKj9PD2O/j5CWvuIogA+qw3bQGx9io1+3NnaV7
sg3BzwAGkWcBC9xK+pwzqH50UCbPcEq9jZ0gTKhWnloXaqtbe+7pUR/eLt28YBr3NtMokO0ZUlnP
dVTfA2jkfPZDVzqff6v3tuZNBOI96epYPQEyUavjBX3wYZ27nEXh7yqjpHxubCvksZSSlHWCBSTe
4jhJcK9oRyoHEbBe3/WMBkynqfBfuLOYpADuXq/pr/rI4zp/8qpj+r+aW8RlFEZX+qSvDJzn6GFr
8UJRGkdL1ZpPk+mv93nhM7W08iF8kvVLM5QERB54IG5CQCBBC97TFoRgtO2aSqMYKCfwrO2OlszV
GBJuszyYDZjgRIaZHB8l+ylIaA9yedM+CyV8lhQ5Bjn0J99OjgU4QPA2thf7dCM8m0lNAM3GeDTF
KSkRIn5gvDcNaqacyWmWpO0udWIeTrtmpUWiv0+cbGkDOg5EltrZtolSV9zgojvvU0UAKpha5DOH
q0o4heEnZuNtb8Q7fT1nfluGvrOWbuBfzWPgh5AiQdsJceVvUwAXGkiBf/N1yVXWtrt0difTOUxb
E8v1ECQahoHkbPg+x4TZuLA4G4H3yWRrJKmMr5hu0HX1j78RI30L1JSDuP3d/QMGRbazUiMEGJob
iDuSNuF9oIfZE6aCuC3vp7ratKMcxh9wRE3iJUMx6EE6b0nAv+5rjZFALlcQy77vFnMl6an1d3cV
jzjSpGcdtzlC8nuo2yKOmBmqWNS6kk1epspvAIXFh23b611KBkw6Nyl5xFOjOBXc4wAs4o+fM6VR
wJo14ZD8p+HSayUwDUr0ikRA7GtbAqBI18ebCB5bDcNwBRcfwtBXLNR2pco5+vWiQ0mwH9YCalFs
UokwiOu0ngBAaDfhk8tZTU0EobwdMDRRySNL/OfdpIINYarTXdwq7iQa/fQjsQtRzB/pkGu7nVho
u8LkNC4bpKWkGCH5iJKsuT3YGZu9ouA1VMFet5e2/IBQ/+Y+24JT9gHj6jUOHjHLtOAbJGxjpz9Z
lcFJshyybbbi7HL4jKK9a4GgysvuWoEdgeYJfljXvv+HkafFEBd7ECVKdE/R9fBiKvk03tLvMFB+
ak29H1Sx9WZrSHnYtUrubSbep8vaMEzDExZe1UB50FcuRR5TGSzayZ3e13hQtjC4PtMg0hdofFWP
M8SgZCnix67XUuwxhBEnWM7XoSVJQdIUHTfnmcb9emPA7yRiWlmVK0YD4D8++zU9gTxTB5f65yWE
pBxc15G9uOA8Xitzw3T38anKmNfEo1W/7b3Fgr0wa/1vUz2RB4elFitQHAM+o6RPjkwccGi74eGv
undh+KIszb60iGgdVEVo+YkCyrzdgnai4I8pxnto0P6IzKPoD2OZDdx9RgTGCtN6mP01APu1m7Xe
CyijwrvpkCjn3nuKYk5KoGiYygTLuB9t2gRIBHJBncIZMBV80+WWOW/uo7gv2Vy1tf4VNe4OlJHM
tMAoV/QCK0C7yE4kkHKfgXPgkhshhAsAtNm4y5x99aWhebmMjUSVaC8e13pHiovb0KKkJdgTBNWz
MbyMVvY48UDRWnmssDlp0Kq4MYyzo7H5hA70l5SqE0idGBT97rrZGw4wX1dKHfcLBPbd6S4oKJ9q
GYT3MbW9O012p1xfW0/GybdtwgV8Xml8Qfiqy7pfMvZ7ZGQAw+RDaHAZ4a6ItLnBweJqo77toarD
AzS7hzfloeNH0aZWKnVq59VMvYPbq/hb1Lj/BhcZ+4Tc8pFBJpGIMR4Rm8FsJSHYXOQ1g0GWD57r
I9hUpi7+3wsd6bpuzFrQCsU8BTMxyHwRIE8WLkH81HTvy5C35WU/IkmQd+h6h4SB+0OopbkhUP31
N21Bszw9Qet866jMoc+r8JK/bLmtc/W1fMc4u7607Lt3IILHNniTGMRZVKpIM5hlks0hJyCKUBGv
8eQfgLc1O4G0cl0cKbfYv5Hfoj2lZFlUOB7lG0thbJt25nuQmX6FgIvmuzz94wjUQkysfegXmBYq
OxefG0GLhLJXlJvzGEvj+OizULlS/xzOc4ate3cTuN7e8mRNuNrKyZbXbQ4sGFmd4LqivL11L0a6
4jD3NtDcpSe6cPXLMw1K6BD6wLeiMxLNlVnM96k8DYmDaqCez0Lgl9pBhi66GFnWmPMtGuj69vtJ
Afw7m1evFPFXx0M8fw3rcrWza+wjv2LXsRMhOuhQ7k/lBSbWbBvqLZ5v5mdY7tRY2ZTNrTdaP1aJ
GFu2YP4Y8+OCF1woKWxicuaeOGYo8FKTfiNORgfK6ECCMLR0XJlwgn3vCXnswQX6uPjSq5oXYwKt
OL7Fsw6I2cWC9K5pt4uT56jtlhFdMnuosS6GjxLQHt7IDWhZsuFhlwcoDN+TdsSqc4MXL7fol+FU
ftwQKz5zYWqUUV+Ji3MNz1Y6tstVEn/P9nU6nE8sqtgc/j8CgYSSejfDh+jB8P2kD6HCRGR5pCD+
wh3g5Fpzv1Zu5g+Jknlh55ffLdDat6dLwVrhOOa3WjNwCab90TfIY1/RCGxGr6gimrYq2b9N1guR
prgLpjU1QlKXADOu+zr1BjDdv6C7VuFIeczNQqGSiVQwZ9K6HQfjPyFiKD0y1W/4UO984L9399WO
P67HHFs+IXcr/sxXibuKEaeEcRq0nU5fpbXnn1HIFM6+b6OMX5pZF+qehWca+Kw0kHaMXueepOcg
B5UPCABwy5e8FLbz3RrN4W7ZgWp9T5eTDIOeCOtXJFVJEmsL+eSKTScbs+47uxp5kVYoI9XF4T85
xsUOF7OKczBX2PlSHKwnQRc+CIhKJVAVHsFiaYnSEqQoUNtax9/QOZLqBguDHNM3g6GTs5J4EkaT
TFN4u9QmX6ty/ZmoXPk5Cml4TeEPaWrCumbRmdVi99MugeijzXZ5Cka7Z7+3gH3v72/f8zQzvjdq
3RNyJ3ghWIYe2D6FxxaGMicIZUMebAXN+5aoWXOGRVjsdBmgC8/76/Fm4LP4Jma7N9iOI0cMExvr
c6d2idR1H0hcWSLFdRhAPfhb8XxW0ZuqVkGPpfzPt2GR72gGbg+HNyb5C5bjfrn1j54x+mjePOA5
pEhKiOIs3dIYBpN026PauoK6SdMdNKw3wt412G/0dCCjKTyAlbTMB7J5Ydm/XoKYYeGEAik/bwWo
luROlavKsTbOLGPx3cIR4r2OB99WNEsSUVO3kh6hiBJ7+ZnHVQkURYQM/9jkYiqRX78AU0u+mzFo
PzgUkLFc8nkvBhrJsy+QcHm+ye8ohA3kfdECuuZToi4ASbWYIlJQl4nXBOA/jgcf0VMXO//5ucB/
qH0VfwAXfK2vRk8b2zXvNXJ7b9f+9AGsRrIbKawv9WymC8rPCzJp9MPYa19mbInAhN3mSIardCs1
WNYsMvUIrHeCWVql3jl4LfKSnQr7OLdBwj2/y/chR4kL0T1wBmwg/6kz1aVK9wR62o41JvwxLXKI
daM36D3nsVd2D7oCq3HGWisgOC6aWM3y7xLe8aEvrSp54zL8NNHOr8Z1gtT0RN4jxeo5fKFAGvPh
w+sIK1hAP0amjMr7U0P0pdKJByPIhe2UUbk/2qO50JjuCy3M5deOxxhwkZBr6g72UM/dmLjC6oRp
JUOf1wdpR0xB20MnMNC3ikfgThXba0k/rfSGjgd4E4kJKKcmIYaeydfmR1N2cSh9+A1vtZci/ERd
Myq2pT3RL5REo9HLEsVxd64+Ninb1tyQyd7sMeEoDi5qlvaiID2vl46TP8o4k6j2nrM6FR9ot0ix
l6JeFATOnNl1KaBGApxMM0Pyod9KzuX+VECjCcDxBxXLnBWOaBEf6bQ72ZGT/+81HA9G/11DU0vN
sf1D+SkBqUOUHjSGPH2ruznwGiKL1hNzzgVFLrt06BC2lGTzHsRFgCJCD5PZf3PKHfTXTFnCNEK2
TWZ76BqqKYE8PF5TBCoaabRqU7N0zldHcBMMgC2JbLk6BNOA7Wke42CPGtIPbNdNEniw4MkLrxoB
Yn0gclX5eKPzjIuWcBVPcb0qZGgeMVV4GLwH4UkASR76NArCh9+J1kws2ppUPovD24/J5DmBXAM1
Vq/jbluMBIf8fs5DoeaeSEc4JQIs7ca5MPNs5i/JexNIiScsTfEzo/xHjEPdAk0f8fZjIQBFbB7Y
+D/tLK3sLzMitK/Z8i088fKyKatv+EFXt0OmtqCjUrkKjIV78MqRFQetvRdWMZNECvw3VVxwfPcC
/BVN+KgfULi47bRIOL50i2UhFDS27UhpHwDaapNmBbA6khe2bCO/z0YnXOEld2GkpbGS3HRYd4Fl
Oh8Kdh5V01wt+sJnxlP2SWokvdV2R3LH0BoNeVkxDQ8GxDhRUI1MvzTFzkJURZPHiyUVracBK5bq
3g3dAynRDULGS1VLwc1nAjPrNFxuixyICfGZBIzkayctUesQQBZ3+DBFBarwlU5XDYB+tX0eVwqm
XCXM9NKSJEwnPtl0wzRBR156T6LTI2K23KSH6wtKFZBvrdJUqAs1TrlAFZeScYgyw8JKcROwyw2N
Q25v5ahpeBgj14umY3vGOG+imEodzBWqpbJZauIZkxPWDMz3ovSIlSBjaGiYdvKNO/+P3iWEiCk4
+bePxQbtbm0czpoN+R9ENCP4jPycQ86rTa2+PCsJESrttrGPrPGcNRjCOLzp9U51ifZZStESQUB1
Yl0nfkBbkZd22VUagN5uMnOkfBk7Q/1rrfKyXMLcyiaktCc5XbXhMtZNkm5aEnolTEDaUD2I6qY2
ndatz8RVRvJ9XNSpFTYIWuUVvcRcTRH3m5nt92Ux2xM+5i6LkGc+mzKrsZA52BvHuRe1wj50PYZN
5M0V60sA5XL4HW5hDKNDIKF8EnJNrs6ybelCO0g0uLu/DxOAQ/Q1jZ3PpPnWTVI5V457Ror3wB7L
YnnygRgJTawxreu8AEYzojI4Tbutaw4vzsKYqO/M/Ox/yL0PJ90Wgj96gyKRM5d+fYBGE/4ZZdkL
k+MPDLUJYqGqzBIeZmjfs6u+qcvj/DIiO6GiW3mv7nVaXr4L29w5AH8ASZA4MzWgVfDjpsPACeT0
UbiA3MynPUIH4e90FoenS1CoZ0ofREi6UA4rCtNubgTWNKBeZMgjTsqZByvDNwusljvpYL3wNoNx
D0Fr/5JjlAze6NrzPiuSwYARp7+Drlh2X1IbeS2Qh19R8alaBOOeuitJRm2hYmkxsXKcLDQvFcHQ
9sJnjyT2YfjtnXeAgxhFM9AggDPUzJHZ0aV3yIIeXaj/BC/kaU43pG2lpUX/EWEcgwBqk1atq1Vm
5Ck6koD1/27o2kWY37ku1YmO3le7/6W4REMssryKthEF/4yaWlGpPzpn4uUGuRcWJuN/dGxXNYcg
0hpsNPw1aBHdvMuQez1BE3hfH1Ss9LNaKkO2MIb96useRUEn3S9xTvcrUsuw3fAzhmQ8Nx8eAScF
AeBYrrDh7jpvv3H9fFkp9VOLc2c0RJjRQRDDiiy0WtXgnQYQM4AWUFx3gFaPWAczevEISBI0d0LB
ieI50JjGBYbERExGklhLusC+8vKifgm8ZjOZXWIsHP136WyBneGr90wT8TWnY8oGV/vk/ygLS/zJ
henoE2IZSf+0vo5pWlpUmjX7z0hC76Mnfq6DxsgX58bsQrZ6xsa7jjjUOWq7JsWl5IFi+EyS/75n
gu+T/eMBCQiRqnwR02DImbn6TZi8Da5wwz61PkLrRh1ANqrcYAGz9dC9HZiM0xUc+cN25RsfE8T3
t2ohdxbmgYC8dtzb1tvUYdsVDOjXK7hGil106fFrq05VgCKYFJcYNNvIqs9ILuFNTlwi3JfNb9BR
GT2vvPfH0Zqe8PlnD8ovwY0dnBGmjmSfxgS1DWWpZJQhiC70jR3VUupjrT4U7ood9sknMjDVwXaI
2NU6L1+hhn7AtXIr2bGJdXwgPUD6ZKn28gK0WB44C4jhTe+l59lP4+3NaAtk6yWFCRF/O4Bm7Fao
6Qmte74DB9vs7s3Jxh9cP8XiAheXASZlWny85PWVhEeP22kgnQi00ARXt/9y01VorgvGMoe0OR5j
StOAdxvT66Kq3JtcMa5JPfXCIbPP7s28Qba8lWcscXmkMCyfs2ccWMhTQiiQ1+dafgm1WF7U9l5t
/dK9cCtini7b8tDr2wN1/Fs680klzrbghPeG1TPBX8KfG3dGouYseK+RIQv3KBiUBC6gy0oftNfH
//U/RJrN29qxjeAnev4K9ea+5kUzvG5GqZA/QKcC0Pi5KNaQcDzaL3nvcOKkghApf9zYrOa+6juT
MbMqBWnmr+gxNxLrRjZS54sbEi3NMk2/Pp9vDBeeu6ik5SZiKbiCKctMwYi1gm6TqHCU2Pr9QCbv
gQ/Vbr/7gNA6DVHq92tSN40uXpmmOQE28xG3c6m8746JfoDvPJp2Hsq2qdycHaG00v/kZ6/A04AM
9KzkHh9XMydwfvCervP4c2yhQhlUOjNy7HpCWLkuyIT5eXvVuYPHDm3d3ctYJoQ1vnz2OQ7s93/B
486GdfY/tVzhAAJb61pzZSoYsC3eUuzZy5tawjDTU8jjIHAkYUcSaA2la/OK6LCayqcsJVVp+4Cf
BinCIAC6yZzKHanT6dgHnfJ7ollDK5muT18CT24tTCcnXF2n9IT1Rc5gXd5YLdqSmtGbmEHbvmBl
YBmdlnzCG7PQta18W4zpr21L7EXjiyOMD75lOfBl6WDJCQvnBiyikgXgTAe4WQ6ff/4CHIqx2PEQ
ydwhdf8bCC2G3z2hZyZiaN7PADYc3nayyAqu7Uw10Ixzw3DfDWbLdc5EufsUqzNCb6KBDVgN9XXU
9DjWMMtel0Oa0/6oCMKw44MigooOn009rgy84RURUo2FSpP1RNoL/ut1erJM0kKGWj17DEyhxbpP
O4xxIMLw1/UsWsbWdnYuieS+RPQoh2ySl54x2ntgcjD2NemWHzfF18u9OI87bYWaA8sG/t+DTF6o
FAF+9pexWrr1HF+//HVxh50xGEuITPe/9ul5Ec0KzoemBRZRNrABYhkxVNnc8/6oxRlH+UnvGyI7
f5JkPc71QFdiZpANEAOzNd/J/0Q7REsE+2i4OKOLyIOZsrT05OGbKvucyMO6EFZPJe86xGjCFWOs
TEpLfvuX4kKhMutKoV8hcO3I03Yey21rQHhVylZ5wEnUlqYTl0RApEZTmIpZEubL7Y3q7YAIwq3W
jwpOe+WFZQ7oDBq4z8fqwHEffC4OAWUiegv/e89/xMATHbX3g9XLIGJ5kujwKCaZ4Yo48eweSZH1
h2p3CYPY7UQew1ARx2YyQV/rzi19efJsfgu4dqTDW5Ym9sFZF6Es6gqA9hvoFgKcWpWD+dM1Dicf
76KO068iXATZ3r02kp6QCQV138WOZTFY/g7o/5g9Mn1qk7y2qJZweYs88BK4OcXcIohZN3f5m/vV
FWR32hBxTeso/NuZy5P7xjJ95QX27xJBOlqrE/wjhbmV2bX+VqLovyFXkseZk+VTrAhk4Bws5uAv
ivVZGHLCsl4NFH4N+3R4Tj4y6fYdGBCMiWGtSZVzPnlgkC4Wy5stApgYBpBBEQwmr2Rzb2hsXpFC
1Apcqf5JlLLgAUoWwmtGAjzvrNEow1Q7j0W0tK1xB943RNnHuvNIPLEdXwPfsgoQN43/MwRYR/5V
RS4st9W4ASL93xxTw6pByz3vl6fBawmA8jmo23x2mZJt8SMbjvLIE7VUMhcOnv9lMcJknzffVpc/
3CxzxOsGJymKDGhak2Cs21Xut8LAzCu42NsfGp/S5SOoIsCxoWw53vFT7wDuztCgXtMX7dk06R0B
VKq6c31V1Xmb2kXsjS7aDMVQH+NN2H0noZPtUxYqi9P1sGMNtungk6FX+8tDiOIajk2xzl9lfqEZ
VviHWhSttQB1C4FwzGfbaKmNIrzJ0mx+LO1Dd/eSkUe7bZHEW7rG/TFb6V1gE0N0fACSfGUqdrfL
OzMGw7uNe4Kbv/ZzXLrYWfhmvUiq5N0tPwahfagYXiu20pRZw/lPlbg/gWOD+a8U40lvi8lWS68x
egcNp9SewcA0xspMcLyFiDPLkKsaFydyJP+VYCOLgT+u/vyTm1OuJISE+j6MlgSitA1Wbkqe1Sm2
Rhdi9o4ak5tofas0IFl5PF33k92E9mz3VXoQdQnQIg/ak6yLE7OhZFz1PHLO4tx/tY8QGZJ5Ejs/
rCW+ykSYxoxSubsAVyZEBOAM5IVzjVztB2uQUqzPbVjG7pEBXprtCjIyEXNjJXzZSZ8VPzPChFbB
cb6kjVrNhwlMJtbAICoRsTktnNR9dfJDAMLuRHXZYX7SRzRhth1bPur24eC1506M4WA4rOsCst6+
rUx88SD0Lecn69Mc/rd7/c0wQg8x8+8akaXdfoetg2EEWuhAsq7AXFg02Z1zMozMmz9alCSp2kjs
L1p/d2UnFMwie060fyV284vwK4+9Psn/BG9DnLVNcyO0XeFnBfqHVYb7Jn5mhhH57UhMtRZ0Np9k
WopIt06G3RPGvno7Um8THN6Y+tUmw+oRXtZc/1xxsoGbbf+Rx9hmDKq5fypv/l0gQV3azIFa32GP
sXqOKGWpmOR+3m3seVLGz9IUo/QHBSa5NjnUmHBx01cJdI7TH8YGJ8h/HlJPWqVt0k6O8oPPt4Cw
NHAdudhasPJYD8k4uSVT2HEsVy7Rm1HRNkXWt7w5gxDW+B5EANWfswskpgm4yJSwmg4LG2wt5fMA
GkSeo7/m7O3o8CiZd4E0gkmMwMU9bLaroMSFzBWryNGhq48fG1mnHFJB9zm//KYQJ4SWFKq2h2Q7
pk8pfJBfPc056QsAkQeqcYOI7d13rPYgF9Fylht/VEuPIdswdnBeAI3J9GEgMWigX982Soj49iMc
p5kmqr61OE/LdFeFSzYGs8OfoJOjtl0jYZNXcWHhavFsiSTf1kag9V1SBnfusfvGOq4BXbZauei+
9fbYhU5Qe4URtpefjIwrCq0TlkEAQR0adfBQ8TBDYHwZiKbR+HiQ/tq4l/azc/T4gARKC5SLRn/k
wGoqcpzKkJvWCBMs6vMtyae76IVF/rsvpDfdcII0kMyYjQUcSVcDMK3TYqY5m4Pf5jwU3DNv0GdP
f4FcJt72EuQ1d34FIrjK4J+TVhBBpeeyIEvaIQTqJE9G+X/O4BWD3spWwwJj4+qaTe98IvARLsik
T0peC7jvsyyVDaQKvSQBhQ9ytOi1pt88rzAGJX30E4EXZVNJorpPqOb6Uu+AUQ7WxzdWDyhYe4z/
satSSJHuUrAHFgVxFLAjzDVIoDA0fQfbp+tpLog8Xanpp7/IFPQxjAT4/ZVPCPbK/DSdCDIyO1PN
gdWr7+WTfChlcGTsAvGcHXME7X6IwZZA5PmdICbJnDIy+Tz6klDqIieCmNoX5gCoWgaoNVKf8EG6
8pOtBquxloMFXkYVH9flkQ9LYWcdD4htIX8P+/e3mkDhKksbnL4BDpizRSAv0By1eiw8WlDgsRQG
tu/MczJusEyIR5WQdz4ZNOWAkGovZKz6S8y7XnDbGrpttREHQJug4om6JNpvxDYwlR/1WDjSIzwE
/fJoGjlQgRsXkM0XU3KU3CbWPw41o2Jl1iSl0Kwj0pEkQvpQIy68hKUiJLt7Vk5XDS8Umw9DClG/
0MwWssM4e0+Z72lamzNl6+0TGecCQgM6qWuRMUii3jXont0mChZvd4ypDYlP2cMq7oLSFxoMbWC0
bjOc1x3zwHWIkfjPsHyVVq9iNbyLZ0HubbgXAe7uqStM63APug9i86LkYejsOFChHxTkc2DTVD+8
dm89VJrGX0efzc71E4QRsQYsOpXPYKV+shqegpsF6AhbkCTcm7VXFjX6+n50nxmYizJd8crM5Tpx
alxXu2GCIWxOb1h6psIfHCwH5BE2RIjrL3M8GKsWKEFIw/mLxb9QLHYtgjKRanrzkm7MJntGaHC5
KJ1luI8MWuh/AEiQ81bvrEQnlADkVlPPtPVUbnmrjCe1PJrQWrkfUsMWK33c6h2Pk8I8UDMeveCd
7fzVCVk5S6g0dGMNSYasXxYjD3cr6n71jfd762XlluW41VEoZPHqX74bfSQzBw+RusNqBeyhmuFz
XbonIwm5w6Jl/2zNF8syfi+HsNB6FdvhHrrYX3h/YsubfwbJIcyQxY/xCJOGdQum+Js4n9pTDup1
KKndv/TD7nmarwHPOz62kgAPDCHQWel5B7CduipUM3BROgGvYKhev0kjwVmqCOm1rkiDfTJHpnjK
kqx+vuiGKfGX7WWbsJx70NiJ6KT7Yr7ix4pqFP7NOpaMRuHFkassYEXGIvzzgmeSuzh2eYEE3Qmu
BYBVHiABLkcchO+Gwi5jVFillQAQBAevSSzliqQGphxcD6zR82lgl+6Q5NCgF2qNWGffGE0Blz5u
Sd2XGqzrVfKMXL2DekZbweJo68CoKrgjsLlB6Yq+MuYlF/u7aGl+VSJLWMq6EUpuR610xDqsCYM1
UCTg5VUyoZJB3EjmpzQhjntziyTXsPv+i+q/JIXISd8WCBRgiCL+uPV4XVCKtgKCA+bSLoTkqUdn
N9Q35SEbxzvnzF5n5DcqBS8m54vxBnZYaOx/GbKnboJwXcXddmLgwXds/f0NAzvVOdZOKTdBz/14
lQzT5KKZpeDf8VGfOkw4oMpkJgb3nC3It9zRLSabQSjw1dVcj868kO/hH7vRSXq+SqFlK5FoHFXM
jIY4N+XvffcINa60X58MHSQo5Se8u7W96Vye/zdD4B1fjRgfZRS/2xkRBfIIbtCxWEenrV4aYBxu
wHAqzNNsLTrgPdLBMxhW9b8gdV164hcbDjrnAv0yZx4KhiEim2PUBFAPRJLF5cFTMZ+Qh6nbTWeV
ajYXjPmLYzWoJhmbGduz8kqLBVJQJgxReC6bDAaNUHyFVdnFaGrFgUQ0nrksIewEv+zZHnn00AJo
c+Pl4AdqCpUw3a7EUsb/AxQR2/EYJcz6+rMCwZcsGdLjIm7Y6ovRAy6uDi+4Ju5eARFlKwFO9W73
7APOJ1ET37y/qND97CHmn6DGDwuxjYoMiM31ylxocIzu7PCK4FNpBtLKwEMf7s4PT39u5avcqFc8
+UTRqNCeYbKaTsfcK4wopF7dcbUWAimNuexLYv/2Zm8aG9YRSmj5/SvC97xtL1aGWq8LsTWBVNMn
AY5Xl0F2Z8xcnleCYEVWD7zNcoUQXTJ6D3tyGc8fv+d4Mlweul9/lm3gCbYajk1BiuJ67T0xWozQ
bdd75gimhgldCjq9uZIKtkw6pMOCUMgrmvjL6RFz3RK9EwLx8fL1+PfoiZcvFd82PLU26EWo9luc
2dvLlCfAoxYg5M288l0VqxCR9jrrliLWIBNzcJ14WEpXoE77rWHi2rk9dii5NgE9oF8MDMK/aNqt
iyYkHE1KxkrIGlmVD36qpcKhR2N/cAQ7LWNiRYtuXDMoMthbJwJjU1OFMCQkwT2YbiuU2zNlAjSC
vS2sT6436Pz34g3sbnEVQ7bRdIn1uga6Q1zuh6F6SeBM2m/qSpQIeYgKSHagXZaVlTCcayzkGAWi
T4FXWjy5H8abyBT4lWskQ3GgTtxX/N0UEU96Mu1QYXYI5qK9ZhZha2MW+EIGB/zNaZjVQ20scYDI
lICmJQ6iMwxv+x0YNk6jxsc+TddLqV+K8Krr0QCzgKpvhsAU6TSQ5rxVImuEk48ZSfVxDGZxM7N5
0s1Hy9aH43n9aOpbPtrJkMdXLLU0ST/jMAWs/dItSFky/P/4knU5BNMG6GPrmbwao1uG2ydIxxwR
tQk+eX4K08vRt9L+weQ/Ln7MaqlGB+KGa3U/LNfWaD+DwaJIuN4nV0uapPp/tYLoy8Im69Ad0tZE
ptd3StuiN0b+spELUN4yDF5dCQ0nH7JvS/irDdaTnCBTRduyKD1UZW2yPl2OxVnns17OQoUgC1u4
gJXfvmCO4/ZuXqysMNTl4upco4oCZKHBBGKLatusBMsuRvYeCocrCrxTilAj7xM9/80vMKUTTeik
oQ+7VmNaTovygrBg0lmX+U4kjgxR0u5p8H8bt5zDHLPd/4eHs/EbbwC6+bYIiwOUZlZuhYO+Tccb
sKCHqPP13HdVBXasuVG13Zbx2ZPTsBzIdwgYDmFYO6aWJ1sautaL6Xk/lv9YYkX2ac8E6IN4MQqF
EMZL6dw/aOW8KP+XPMuxJXRp7QWSODyX6fABxCo4c+NChbrLmyNZjuOQ3Rf8T5Waj2R9WL5qYRxS
Q09JTDZ2X0n2i7v/9tdH27emyrqBKnneUJ5lnU/3QcsVyq/RAUciX7PSU5HuicIZtgzkEBrPehS5
gua3cXOz4u8jlqGV0z2giLeLc6Ls/p/ey7sSaS0z5hzSv46cgntHap7JAM4rQ5TdUHhDwGMIGy/V
TY/g52zcO+RG0leEIXxQPuqwrW3LnW39unPqBTdrC87VXdKZMa/bscwEAO34UWlR4rmp9cDDFQOs
gjLhw2jtZRDDWRgPlCQoapDhVzz+7zeZPT7kGJtPPWMMrDWrmgEV9JooT2VxgG9Bkh5oBPZoRSeP
HVgkNMuUqSWap+2GN4YcEbKcpsy2Mp7OJAgtKUrVmi7dZoFBPuFBjvEwF4f2O4/04RF5fcz/YE3z
DckpnKBw5oOJoEI9Zi6ZJSx3Lvfau3eSKSGSsK4IdUJWv59mU3cLuvAvh9q/hxbkAX2Qd/s5TAsZ
rsTgE2NTXfLdWL2zo4KtiQV1g/koqpUNKwehG8I7cfBs8MVVol+8e6hgawiPHwgSUqID54lu3+8i
nQJRMKDfnycdb2oyVzywDnrIRCxv13AEY0dp9EeVU986UDuTx82aHixksXfXEJfn9+lyTmfovFBy
zx8qU5tC12pViujrlFWbzrtjcKW2ZwgIP1+iu9XZZXaQMwDApXAFuEKna5Ia5VxlSpACOOZ5Tqxk
jPkUOa186fmFKEBQligGVlGhp1Pcb5koG7W8gO3V4OQfbKWE7VXMPrm5LhcLLxM8HaJC2Jism4Vs
v6RBWytLK4k/1zdxMS8A7M0+bj3htkVehBFU1yo56Oyl9TalFLlnMBFRi6vSYqabal83AGWW4RLc
EensS3EYO4X42pJM4A2juVXCF3J64SJAozbQR0SxNQy2c/Xvmc6jFipFf71BTQzAQEsS57cqPQN0
282C5Gu2CygNoTsOJBr0xSjy9xTmyTxPe+j2T3dcZQhFXcO8/yXvxckru8K944lRQPLCoueMQeND
hwVS0dSXZAhDeEjPUVEeXkcksjgyzGgG3yqavuP1BLbjicAW8cbI4bh0RX8cgfFmTkpEoG7kzBqv
13mTfkKqsE0p1VxkgGw++1//8YvAemxILb75o8PjY0chYzNsBZUEjTXhb+oYykRp8+m6YtZFbmIv
NpvXSVBYNAtrLsbvHIBppqnLAJySsGrp/BoJr4yCX0BvbVC3bFU5gvCuIgtpGbr/IS7thuRvObr4
wVCCePGwPRSPTqsqK3BXYFdLNaniWMPaVnc4/w9Y7ZtLdxOwZJrBdd+UJxlJRkPlJuc80lZyVg35
ohIz5sHE+wi02CIxBTVnx1c7mE4G6UnQCcLSmL3yTOLUnCTFfLwENP85vDrhsbwk/zVeEleEP8/N
BtjYYAaemW74PJEWOmDQgkDpeP4Kgjacrim8a0iGEzpAUPtpKpDjIqk3OpCDlrHVYBe6p8nBME3F
5cczvW4lpvNKZRXDG575qit8YbV0T7odTU7ig0oLj4iP9dIKrkVw44toLPqN5SKCi6lj40mWV+17
haMnPi+zqlwlhW2UzYIf9rApXgDVr3ixXN44i802DsXBfQQlVOM2OT6mTwYNuaibHZCRMpOmBLwp
t0ZYEHnlSwXXrqfqxUaiF6a3RH+P1to5ouneGk67S4Liy1knJgkwUdKwi/jn6RCvqKtaisbqDv+R
oW033qRb+SFSrSc0ex92yrYmGC0j5kYUnF4D/mq0iGt56OyoWbIBWoSMhiGqpo6A9puMToAjoX1w
e464oeZYt/hN6n7SBpFvTZwmhQ9arw/RBgLTlqdoJzTygLfH+WIM54h3bTP/zf34zZpHSsfyJc0f
xIRafXkDDldSE6Cg0LMQ70AoyS1FVyqonW6he6IiXtBgUT0jpvQ60F/Fi+3WBqdJlpT0n8CXHOVU
RONkDyDbnQm0QRWQhSK8seiBCf+jpZnoNlrAJYvO6/INaKRyKjG+tQW0cpBVrEtWsyd3Ihbr4hii
MdjGo6yHWcbWQs/EUMvWjQKBwvYBPZV2AoOqyjq3lphnBvAwztLGVsrvpKpnmEtU1bta47rYHgV/
QXnw4NYHk8fdIPmCbQWpYI5bOjnfJXLuwX9Dqumj44Lmo45v7MyAwhwjTm/4HLM7/WEbHpCmkRn2
r2fnvSJfgE1T1hqGaP+rYKw5ZPnr/1LQiytTBgBKY6PQpsRwnA01nw+zwD4voFIfFuWl7WXYm3fG
MWKwSEH3VL5ZPS/ARfl8DenbxLPFKln/hF+TYZqRYpapq5Ip7tQxYwdj3Va1Ma2gJ4WYbrvl9j0U
mw5YntA6MXCpFediRk9jTW6pnQtb2Fdn/xHJhfJcerLwVn0+BYpwGQ6cVXapIZUrxPmiTbypWxzY
VoHgkC+xDEWLHxXT7HYid61APj3VtaRGAOolv3WUXbBTlK8ZX1l44H6h2o9EXK9PLkKANzj5n64T
LW/msB5LPREhNH82GNf7ZxctVjhiniXVkgZXxKvnuTIuIWtK2Ff+YA43iCmY1MFlCennp7ezy3rt
qVfnV6SRhipqezDs29q//ZTm23YbgHagQlMxP/lVB8JOleFbFeadixmr2YcLeZ+Gxb0ftVo//ssB
mRRX5LOyhMHPnJ9zt1Z9rBSMYKXS+P5R8izi6uxxik6HzHkwKgYPZAUg9hPe/ogzZbSWaJpUR+pG
jPAzjpOt4WBWJyUChGSXtjRPJv7F8Pmvk6+bUBbU57iRDAe79w3A22uIe0xYg3ktara3QufJvist
n7YMJ2M8bxUYZ7IjH54Fh6L2cfCMEri5/qtRNu/c0unWEV6z6UlsSHTEw7PLEsjE5vo6k5WXQ/L8
/8QGUhZ6kB4n+bedjAlqdECfZM7vd8aqsYDvwuvGPVOz2I1BmSGFy6S4AwV2lsUIQh+kEig0Llok
siPKp8J3LLtjmbR1UEWZgECKwzFrdC34/dZrv/3oUzxkFv3K0WzPVm/195IQqGHE32VCyQe9+tvh
XTVjGXx+v2IBGHLzvIS8L1YR+l3e4DhJtlOTlqY6H4SLmRd6Ge87VH/yTqT+BB5SPZxT9Iz3jSTw
PAVygVq1tdoJmvGFje4kM0R5ojG24UzDZvDWyZU/N9XexHD/EMLJXoBrSxxIAouzJNlmtkl61VVQ
DTXawEfb5MLB6wjzwCNHSkc0g7XokQS2ze5DpRv6NO4ye9TwfGGuKNjXbWObbnRuwS6VISuLdYEp
3JHEM6tmLbknNkjn+v+TwNpdiiAW5b19FGCadKtUiAHrMSMjiLTZcYlakAyy0rQ5zZTHXBcXSVxo
VKCZSfcrGhUMRm2B9GWtibSBgd2I87BzRvA0eDfp3xpWkvA3gPFdBTYX9Yl9qxI2jwW5NbAoq4Ap
PW0nNfcPxZK1XkZskm3QPpf1/oAx7kGYpxmw2uGE9B44dbl85GhjeKja1pB941unSlm+ydVpdwIj
7jiZGZuzvAN0VTL/600gE4RjGXe8ZJb2thOQUkYqQyngBNp26J7yjlL7Yy3AlUqSiORmke7HIxBO
un3V5voEPtXHKe/90LfiAx71qQ+bp8+FDu7K1tdJg5VkJx9TwUXk/rUsOe3MU5to3sShHjMy2IK0
a/6bISLMAo85QhYv27QKyxmrUrzJze98/Ehdrgk4ue3NfF2E8bUYt98ayISq5+JynQzaiKfBCWjp
UqxeceX9lPcWrfjnDGJey7PdgKSmlubci6FPGcDbNoJooMEXi/WmF5VGgqrIZoYioc/8vVXVmZej
SVwLfEdmhogRcifN6flMCTnuyf16seDAh9Qt0dXFnVTWZ445p2kah5DNB0Yyt02kZlkT6wzOhTds
qgiIIsbRrPSDrgN6eOUPWSVgkNYGWnaDbFUkezoOLGMZTSWOmNivZ2FGPZjGnQi9Vk5PWSv6UrjQ
0qPDXxh+3dK9U5TCXZUgRq7fTSCS2dlBJgLoP8YDg5jTXiI76A98NMDAmYpddYuGARz+i2UmU2wL
h/zwipLmXNAV8ev1BgPihLDwKF6QtS/rpgDXfu437vSclK27rrB0LUirvNBQATspYkeoN6pAzCpr
VMaQ851+WP+hxx8yXJI785dEZ+OeRyJ46y837UrecLaH2wILeq7uYDA4KcM/RPGeNtJiqTN3/Rm2
AWfMQQ0ITRzBdoY0IFKrZHvFM/g05oZkZiKWgjHWdetnu8gev48NPF3EYLImlSTs7msiR3qVff/4
1FFCtguJyUZ/+ctO01xt0bIZCZby5wqjgFGjovzISmu5C1mbbwZkLnRwBdZ7OBCaTsrXdII5+EL6
fSRlRZjrpCwOV6FlO+Og8MM0EpYxhQ260kGgn+peLflD8Zti6wxclDLrttlONmp54eEM64aUNuBu
7NaQITDy8v0MyK7HrVH3/6Paet6Slk6t8cudi5B14eYvPsObzR0XC3jpayTt4zy39HLNIx94f4ps
RTegTF75agni5YdUDCRFu+GPkRbtaBBYDeMg21680Xv79IOWeKIKSA7SJXF+dtAwqd1aql4JMJ3n
7COL99mK4wvGXOo7sGy3MykeApPlCIJX+4Sm5w6K1gY2QSsDiO08w5AyeE4/tZADTcGgKqEV+tVg
DpX1wWalxANyReqSSHHUZSH33k64kJBV/dwaln3+apYOyblvmQaeOQWWcXTzn2A+pbrAjhgaoHAy
DOMzAIK0PVSdvyx6SoRGO170FuF5MnmoJrkQ5QZ+9F+nw+3Hg7bD0jyNgURUp1A71arJ+oqSGeMa
ruAsuDW6i/82ACjJE/TKN3XbAVSLuovYsEadYlovTW+lYKlc2YnD9wz79R1ixenFP4gPk4EOd+bA
HdoWZ1WDVK367ZjI0GATBvPRY1V6+MJf1WkjFC3VMMo+7tUTvF2QpLUL9MT/RnaTmkluI8LlUwJD
k+Tdu3Kn5W4hcjQa3XOO+u8Uz57xo/v2j0Xkb+cdgDQRlqz/2wuDsqEq9HpuwU4spMumnhr7vB+9
Uf1s5iDEpcYZo27C4TLgCK3NUiNKxFw7Z+Dgnj4xbHQma3kmvi2ejhVYr7El7jG3kGQQISvsQZ7W
n5bMHq2tWPFcQQBTVhhNWr3fqCDkjCKPkHTVzzpSIlKBQrmtZdfIFWrKK4V6/mZnFD2cP5ZtHmZP
CvrhErVjYGsbuAMObBOFZfSHIYPL6+FtaZZHcy/nx5jCU0kjA6X6KA/jZOVP/XQNoToAoAFg0g3G
xLQy+LgT+2O6pp0Jd19c6hhmAGqOKN6veDCmr7WrCut4yRNVRlH++L7IaPCNLTpc4wRNbtKo7GKb
Xj+sAMDNNDv60rPMKz8rPwFYJ/yf37Mcb511zrjVuT/ZidbGS2Dwq6lC49kZn6Jicf2z3pS367xS
ZVLtZqw4BlBT+fMWBtkaKuhhzrI4tBxaFw33yoCRGolgcTPGp9Mc3SdP19VFMkEFBBGDHCvEjaZ3
6n3RdBklbj0Of8mR2nlmBGbiZAtYg3qDqYn+qE3RfRR/sFmBxfMe6m4Bz0aAFhlZmFfDRJg69nNf
s59TJaTU54gp4YeIhliehufrI0C1oh2pJ/du7V+/7vX/16+MzkRuNW3IGHVUUglTwPuzeLuDlCZg
92q5qfm+bA7PKEGNJLBsExiC37H5849O0EhgUDBDrIb0MW4xpt6qB7QM2oIly7pLqAcnyVjH87ll
SjOfaKSy1Hvl274eJmu8qsILIhl2+hyS1l1G3H1kmyLCPnDePVNa3VY6+9nnAdVw7GB+PXWLEzHY
eIS2/KSZ62F0u8U6Jo93/hiyhvAUQZSgQJaJnB6ubow0I7aw6J+tlSVSDz5QwpdUVqwGu4V4GGPv
4HK2SnTBo6+iUike63ZcsjxdnxpIXgglieqPQf6eHiYjMMt3/og2RMC1iLOq6OLn/kv5ytnjIxRH
ynXpBfIyLN4zmnkm/3p3sWqvOwhSUgne2aZCHiohQoeJHPpy9UIt7ummDOLl5zQS2O52egyoxdMH
tvQ/rW0QIdG2ek3ZBfE0q6N7v7R38tWpVEWAXEDRMJsT8FGxacv55OOguMCNNeLGM9RQKCRI0F2H
Q6uMwiNrEHYK+inae3chbVQYZFBJzlspkcnNx9kqpwNRNM6p8TQng8G1u27qtLgPxi6eWS3NywVF
kvjJtoaWny6m5Qu3LmZfWm/anQ8PQ4YbKG/+uG3RBpwtkNOX7e/vDQHyZG/UaPx18P+gEL5LvEET
ujms/Mp3XdqjqHiOyz1IjcoSCHKqSFN2oq8TjiyDMe8Tt5Y3V2Kt7Jjesi2qQye6F31XNqUHLFQ4
ahshaeghhnmDWGz8vKvvtJGIlsjBZbn73WOZ797Rz+22NqbH9V3uWhpvHf0rV74Lo/4g9hLfbykw
Ipl8klKfTy35tDlwop5eyw0ZYqVnhwnC1VQRsHKWPxO3YELgmmA4UlxDUdXm0rekTlBahmlB4VTv
2EGKC7m8Lyb0fUiF/CTEHV0ZtBwTjAOd8g0Jb3824syZT48zKetWKeDs4paYRLVYe3bP0a2O/7/d
/bNo6ZsruOQcS4MY1FhfJu0jgY9KeUreu6rpMnAX28qt248SQr6BXY/u85D0KQd8JnGBocTPCmpx
3I6KBvvwsorPVe2dtnBcVk10LruTBjXfJbqfdXUNDnH42wS2UXiQGPtQmGhdk3OfI/yXbdwoqRWK
vQyG5ypsqo7UKVv6qTu0Msw1oUlYRuz8CkgOPIB/p8t6eTDcv/wc0xk/CEbfFX6dJBYDtWMun87M
9bBcaUf6oCKABijMA4WE9fug4pK61P9IhgDWen7MhTW6Vv8KPaTp2X7x97Lfg4rU1k3pJnAr7s+Y
6V7jv8BvTEok0GYtgLeAlJf6pEaLzX1XUnTKfgaUT9BTcOScf2IYbTkPEx7aaNnG41F/dSvEHrwC
7fauI68UcFKLIoh6kQOQhwSmCF6AP13fmbhpjLfu0ZsC7KoBCT8z+2ljqaW2IuLv9BPc/XlEoN7f
pFBIO5sc96Ft/6LuWa2KF4M5CYZFNoGVm18pIIWmJitJ+q+weUp7C3r5/OMqSxeWlVhfZuH25gVA
SApnr3AD6x3bly8C9f/YassZclq1HY6VUjqAf3Cnaz7YUTEi8LjxsG865Qo+XN9z+cMW23Mgdm1Q
UKUe5EWkWeIvhNRIUrjtdb2w8ru4Ed5mKusXJacSFXyIq44IAcz6bks966Vher6gJDf8FOjBCYvi
yRTRS4P1RiD4j5PzJjRePLP5dcO4FETwVsuABjBxG/DOXFgqUfkBhyfbVXaocO5qTPSZ6lVVG67B
uJUBZjpGD0RCSyfSSqS2qu3yXefYBch9o/HQKlDnICyxe9G1C3yFSiQUy4FR+1Sbp98zLAJMcKHq
QIBe8jZrxfUole5/1qaDgGmaCj/GNKMobj+Ac5EO6GHImhR/uCkyh8lD0lPyJdZ1OpnjdkbbAdhk
WREjGxZ3vkmRvakKyGbScZdJYUbkwQghtwa5FoxWgxMNE3kxSpMDQm0p6QWQDhbrnCFrqiYiG1Pb
iXxDpnyqb4qFnZaHio7Y/Y862JLklfO8H9lSZa9Rje2CX+XFK7DZ2mjVE5bod1LwTG2Clqpi+w1o
hvKLG5muPNK2gfrtwkEOKEOWcIfre3KFnJPUNhQ/cHGxkz75sorz1byHQlcqsRMU2xusIRHpNzp/
Han1bf5K99Kqc7wowAWUAw/FjlSk78uswvq8odrjI8/ItooY6hl4efBvixLDPl6OtLBD61d35YRt
jo2Z4PG0+Mnv/eimV+8ePGyg5TTc+5njSPnnW26KXr2fPEcve6bOuaCTNx5bE2YXXJxFX5MVvZLu
vVY/H2RRmsHvqmPZMxhvO4zojkljx7gDfVg5J4xg8MOJysQdzeFMhW+wFDduhob5vbCvN3YcclJM
ePN62mZntCdGF0uiMqIHZZjhyZV04qKMyJ7KiUnz39Rir2DNO8Kb3cGAHPrXtPUr8cqaTby7+sQo
Cu4E5C3qIgyZAKJioy241jANOJ28JA13s5IWa4LJCvFsGwhYBOEfejbxKZEOHjhUZjs9e67x9TPa
sZPxV/f+zi+BTwIbIuSQ9bfR3bmvYkalukdeUwwKfoGxySrLtbADkapVqXNI0aVG9i/dqbMLXLbX
RIZFcbBVgIoe/POfvfJ6aUEVay3uMAYU83cI6a+yy7A6CLvFxFEW9Z8LtA6PeizEWtMueZDfcSoW
ej6GopaDAwx/m9vv0Z6m8HTTuYRZW2Ieyd5hPplM6EReivQh2t/CsGdMC2t5zeud0KsNeEYUniem
zleOygR37XDxly54UxpMZo8zsodIy758L3hzUGU9Z62Rc5hfTlc4PONCaQiFxGm0S/hRYfZmwB6Y
0HKp42zyaDnOr0+ZT0Po4SDSnq9V6KybIzbhM+wG66OrOT6MG2Zg5+CDzrIJGfN6GK23rTEeShCI
aTqefpc5vtlTjC0CO5f5LG1YblRaIPIZ7I6bopo3zmnYGpTjVQ424juRnu8SpRN8yy0yU2sGrRU+
PK0W9Y63yMzbKLUpSl28gAO4JR3qV5tLZJh+/LNaDu8Xj/cQyEsedi9Khd8lSTyIZQ7vt1NRXbnV
YYQC8GeEN6ZZPNSOemccud7+2pktMeJ462trDkWzFIyPSxM0WcFxurvrbx4z4MnuXpRcAzfLi67d
mnH4DI6Esx/ycqBpaF4MU0C2iGRUGgcAYcO64k01aVTTdxDoRF+aCnVpjUQECzGnm1BaGoF8+XaY
A/xbnLvPpm5V3VjtZt8v+kLLuYwKcSHtfteh0G6Fg8DuIOaNZKKdVien1LTHe7F4b4XNWPCUWv8e
A4DypkSpDW/V2pJrQZ7OdkXCpfC9He24vYgk/U5pCZ9BrVOrPzGmxADCV74WWjAkqB+BeyZ9HJm8
SEWpchln8ZvYYTdMZJ3CRYZ1+LCo67oLaWrbLhdVFgQDe1fpzArXzJn9bkHQ4DPjmZbDr5Ddmptr
YxBITdyHDj/ehWQ8QRbyzDKJ+NGG+IG2NjAzCdc7EyH7PI3kwgYfQs9ezI6xmgl7rlIZQIuw12R0
BhRanGIKBLebfLleVpQjgKTfVFqScTX5sArdsrOGRj7YAbw9dnFBW33ETgQBtV2aN7hb3ScrcMRa
O59vEV4oAazUYAnYpcKQpYdKYWFt+H527dRXX6gwaIYrtqSR+UqIwr5l3MEQc2v2IWgl2+rlV31D
Jb218+0WIOymsroGfsxQGBOX+NpBxeqghENAYJKs9kmjvsL03wmQmAuwdSVywIlTmywhglRV2pEN
bKK7NI/L/vjptmM4yP2G9QBUmafL9oWD5mO0k5xzYaXCYwdAu7jXA8CbGC9COLRlOfSGkiZh5/es
S7L9mOOpQPOoyxEdNDbuOM+v34wlHHZOkMIAsDBYy7T3Nv0pXkb8Yq+TZYZaj9HtOVMCYZLlOBlH
7fHmPvGEysKrdj9Kz2kWBClilW46232pUuP925ztsF+t21uBzm7XxIaqK1B3keIR9s6HlJK09sOh
TpO10FrjvNFH3bxqNXv3OYQnNclzZju10DrhQ6F85/0UjQAzQju8yZWw/rB3lZPOrFSS86Uyz+P7
Uy4LpWOmmGElA/SR4qzMEoOTTbBAuvMr8iDJuOwmjE/JX6HDNYkso/gDN8WDNTq82HL9DgZavOij
Rhh+MzPc/IiVCA2XauHcjQG3QELsDUAx2XEUjbUgBFi7o6R3LvHJxMd+MEyf3J3A7CahLFfXdz6F
UjJqPJUhgAXok1h4qaxWCpO6z+hTA8YXMUfdcLrd+cL/vPHvXIXEA7+itnXF6gqDZ6/eUQYVPMZH
e3JZ/jxf6BDQ6jlF7nOSd14lnzyImYQMTePv0Qu5w8KgvErEZs3q4azazCt7jpkknaiY7KQUpXT9
Id4DCqVCcMkKmiNnlJxr+Az2wYclBFKbLSy2ziry9qeiEmo71EN8PH7ctG9BFQXRE7Y1VJth712Q
MiHbFkzzGKEq3TIGNDgDHZjJMlQu5Y4wFwnNOJFZjxvsXvBrvIm/8v6oQFUFbGCN+xPreA5hh2X9
EtWHpoZj8m0mRa2eHS/8bsF7zH0jH+a9jbTkr6mcWRSTZU/GqqL8heRCog886qJN+R2hDmZ+GUI7
bhBHXqIpDRHuPAM/JcQYPmxkuaTfJt5AoxWMvUQHUqJqMa2HclRA2GTxBS34QjBF8pCZ7updCoY2
QzMy4zbD/0ztER4J+hirM681G3B8/RBSHzgWhC2OuAeE8ngSEqedc294MJa890PSkGMrz3NO9Ysz
kyEjT5sWC+wymb6NfMCZNYuF9fcpG7F5HugGMPbK33h1jVpFMnZtZtYpICqlk9jVv3bBwKwkmCKQ
ZzEfocg56cn6ZV14EkzKUa+FYpOyDQTUNorcb+/ZwA05tAqkKe9vG5WbBwk2xb8eDlJqFHkT1nQh
axPv6meQN6Fj1BhhyDIaO5GDLpIe2W7aepEwN0EAB31G2zYiDGyTho9b18BK1+XMqCKNGE2clnQ+
MP3jyayCd4OUM/PwRqe0S1IBz91GFjOoUxhyqA6F7JrFDqjfaxq+C9maunNN9TA0w2nAZzInwpj0
bya9mq/iQ2M/pxMirRR2SqDzLBI5t7L0IBCwkcA5ESbpI6xcXOoteDNEtLpQ0TNLzG6rrdE7/EIL
+v8ROjIfTlPPbjJw7LavEJ1IQ0K3epB3V3+KIb5mdtKMp4332PIrfVPzxRSRbV+wn/e89D/RVAYB
h7GKSLAIRwK1z2rHMGSvrk6fw5z0VxRH0Zs3tXJo+NjvOianyl95PnFwDUSQjua+GpWVu5gI3pIj
98kHpgY5LlxkI6SLJPxzORiQhVVO/eso9PxrGp1/ZCdetZy0XLzByOyl9LmM8DDrinuNdaJvnO0W
65cq0BnAvEIfbhTntH56S8tLB1cQFtQT/do+kRiXDhF9Y9SnIjDpCWyjgCno6rstmQFsfgYzw7kV
/rjCx3ZGLXh34oi7bxVB7E1TlnUO+9QmvL3ktvb5k/PuGxXjq21vRAMw6n69u+Y4MJf6BWyeZeNz
T63hCkA4EtUqK9D3IUs7KTJzR8de+rWD3zIWBmbgH4ENHQ3IIkWA5fzSVV4nwzeQ5Q3vfk4MEf96
mQ1WIEAjqxjFtbla5kZFZJPpePlUqnW7OwDAjf2YMNzhwrFH5dlPc5zUppzapD8HazpxKNASWmSd
pzKLA018qPHUSHaCmnk0rjpXDArk31/BieZ/HWh2o5s51bdDiyunL6gHlo+GdqDjAjcLe4sOKmke
7hyQs8luzyssyE1klzCAEgBr50v/tYKTWMuVBUrWJ///6nLK7HlWOsWRJu7ZcJNnPh6N61Y7/3h/
jPBScxq/LpMP1QPt+HcKGjIN6+9/BexCcN76wRCdsqG3JseZ2jck7JgS07BZSDQcd41rFY1A/Qwz
4oOubiFX1nDRbbYH43DJnMuMGbguyrBrdfT4SBIpVnWAUOK21skDBJGX3OYDHrrCIDHcnYgzophQ
KNDkF27YAEygSGLCkM/hEG1v8oWWBpqTdVXZE82BD3+2qPKTaQ97gE/6gB14xRgYBHDkp9hAtddw
dOtSWtggboHNH+ogWeCPqqrmuNJ9qSixKD18cO6dkEM6FlUGQwYITZlqT2AB3bFWwZPWmRRnoiZf
YFKdd+lboE6TAGRWrW1RN8XnWhfQ6D+WBnD1gEaeaoh4Bv9VS1cn5Hl8qZoXl/sALoajFrvCQYNp
Uwj/WBsnwhzlShRxj9RHtkE+GQMxEMaSSECGOr/FkMUpOI4Bb1NesYFE2qwCaNiTdPJeWYoBrJ2J
g51yGW8C4XueiZ8BZkoj3hDRIYYwwO+Ft72ossEOYA9Urp4Guy7RGiD0+dCib2D1iHSj3bR9UVwL
gBArV82opvoPosVkMs8d1hOcEpCVjoHfcXxEzNPSifQG/3oyXMD5FGo5x39yRjjePLTAwhiQoz8j
ydVEEgT3CP5TCJGMFDLpplhoS/9j3tLdG7ux66KkYLC9TjH+V1IbJqdeXER7J/ZW2tqhncO11tB1
130boz8OtdzddDuNlt31eyPawc4e9MsCmaosJKkRcCSo0RP1u5vV8zSc+aP4Ti7mJrW1ik2j2Oi4
cVwbBjvJVfjVuc4hM32boX78Nh6N1b0JyjkSyAqjIj7FOdy6algiGmpV85B3QR6HXmUN3lmUD+Hj
a4beJz9HUdycPv4bu0aNurXS5TXT6kjivGWZ60jVNw0+G8rB5GK7jYMbMswK4f2CW1rUfMX7pKh/
ICOYzwUQ3qjyBMWEXXWD/ccqPvOywnKweB4yc09X+k7+FQi1DNQtmUZJNiTpdiqSoc0EOCbL3O8H
QKjZgV43gCw21GoUxMnliJYPkHoaMDvz9oTc8qK/F8XXY+H9+u4HGIl/Tiup2m3udOTvixSLjw21
sTTULjChBLqmgPRV2l5p+XRy8Wy8Jns7eT5KasLnbcWRFNBg+6F1MejwO1Wula+z5sWxtFkgSk1t
7XyiNrgPjBv/48TgTY3ZKbdIxO63aHVJsLlRMU2bo5D2prXr2+P9xh/s4PUtaFXV2CSJUwDZnPDm
upp6pSCh1rKv12ueSLfiPHXrlofqWkszXWQ1ivnmv7OCvjL+QSqgfuw069wZa9u5NcjjdiJ9c7re
BQjTEbVH3QrWa1jgujjVcRVYMLJCjUOFS671uaj2SDTECR/SszzBdndbw0EvWcXIt9A3IdX1QC3k
k7562GY2o1DPNeXsGDi0PB+E+c/zOqTA68qqnbF40XXwvHGHj+BVSzz0YbFnSKY4D+F9PuewWi1Z
u2qx6xgl0p/f85Vtdb5O6SrTAe41eUB0AA5CFRCFKtHJzLE/8XGdOp/3ZxyyUrY4ancP1PnXL1hX
8pGJaIMZMoblMliSyUbiH33FTRgNRiisRnoeJ7FEr86vTyOC585aVs9L/K+AM414tDDWKbaGkgAS
se0p1Gr1OeU4+Wdc1cLOPj7K4vLAr7Ej7OZvTnVwJC4UchioJ2gdrX6emsoJQ6zYzzAS5l0aInX9
FHKYs0/s5VxuObijFwVxCYc2GbpdW5/MqOD0X/Z46EUzamnQIAZpgSYNwmxZYjlJG0GTbP9fF41P
tT9zu7PcEbKeFte+WnJlyGZ4pbvreSDnUn/bG8YhbgDGcBKx1g1dygT1FfLAfHBbvw5No8ckSZyE
ZmxvMg29tg/zaTrPPm59NoITRzK1KH/31bJwCOLeZaf6+Z4756XpRlB+ZyQxVUg4S0ULegEjsVu2
kFLJCUJnnDTNe59hhdO7ZdfRGsRnexianmniRxpK7eud+v3YXnGx7Bn0BphPR5ojn16mBKqWN79E
qKDJOGOe6DqYyp7/xnRJEnB33RV6tjKzfonDQTBwQtLjluKGtEnoevFk5pqQHskDNdpJB+ZzU6/n
uLxOqusiqsirFF/jYxFLB5/AFUGlh18jGGXcunjJm2NOZ4dkD25vjk4CbnnbC8Sc/uGfXE4BnaHZ
+EVWRqpJmrw8RfmAjW+7hC5Yt7i4GgVCseR9BrgWPfmxVJemodlQYlWlwSFwCZv8kk4qu9gZXMYh
btPWdmA6RFhQIakt6IHnInFjxk/6erQC24GMupoBp9rP3VRGS8vaiV3j6WUEYX6FVNQ4HjuFgX/7
S4Se7tLd7MTFxivFTBn7Km5a/M8zSE0aqeIkdjGa6300tjKmDZiZE6QsQMF1J76uhZxPBkebZXTU
m0iEw9I7Re9DuL0VdWhXE8oR4EgsRluMZXUXek5BDw6hvoS4sH2Ld4/KK30BwQfYtWDI73dcYOFD
hr91/v0LZwGtpbl6ApLLOXxfw3PxvXLazdQUX0Ttb5AiM/P6GmXHT8U12Q4Htup2b9JuA4Cylmdv
uaQilqf6Z9qfqYqgn5XnExKUfX7rFr+C419L53j0RFqqrcurKk2YH+TfX8ItikQZRzkBY8u/eE3B
ORDIvB0ZklAQfZzH/tivrcYm51cmdlw3B2cT/DcLX9o6BM9WU7t2bg3s7nexLutByVQwFhOdcBtA
WrFsoMtHXxT1CeVHyWTDKOhkufjZpretLHX8PEySGIdoikj4gewyIKIK4sD/skzjph6b+WXY/geO
z25qZNUQnfUudbn6qpXFJ2UCE5Q3i36nNEVL5wERqloqtM2cUNe5CWUAToQm5DwcbG/p0fgY7G1y
w1kjQDssteZUQppXHzo3hT22SfcmRVzCpjoz1SMe5fa2vsdMur+N+NIdFhzs5O5i7jnXS3srk1kw
FRHBl79iIGpkwqcFY2lSquHZLxvOc+XlTVqNdqqhl8YhCE9zF/7ne8KNOewWEApn0vVmidbUMj6C
vY8BP8txxPp8QWySAfzfcpbVtO2E6UeAXWr2MaXWkPx9SLAPpm1KVMIzYnWxJQqKAA/V19oE2E73
GZuzQzUL2ddK0AWfkYRcbqOTaTuoXlS4tNnJ4sjEWYfxXWRI0tDm2yoR/vPuUeKUjQFvLxHatJmk
uiN457NvrhTyK3n0PBeLY383/pcBRglCa3wR8yIraBb27Y6BbccbDJ+Yc+e4Bd63Z5+picWSeTdM
n5/nsyC8FYUux2zbfiz+yhIz7yPUqX/FnM8bzLDsS9hmoUXzUn6SbooIK/nZj+plXBbDTi/KoTWt
iW4+hwWB8KBREzU5JFgdD54VfpeOEHDXGrFY4xd+i5vzl2yGF3HeVrPXc0TBvVJuliJiwXKvAmsM
qMXoTgEn4QFBgkEEzwrm4s+OO7WNN4WqW5XLZP4uidsHesbU3fjI84u9TyDzUPfjczSt+a0mnpfe
hIdwfAyB8FpeqvE9jrEL2hTKOZukMIy4wNKUi7BV4b+abaEQUTtqSSNY/pKatlqn9sl43fLvSDOp
S009uKvN5oLbKZnIsRTZeaN9l5l82qLez3sPGB1cMRUqioBQX6PYE9iiA0rAKiYPS4bIVyLceFRD
uaUqU6wVevonxTsGSy3I+uON3wDSAMyBDhPhWpU3PgygyjdQCvtLnGr+o55nLygtW6IUiM2itREU
oULWDsimIeY5O3+zJcdeJBTLINRPG0yWwUiRNL8TxloYVgiOr1Je6nUSLd5t3CgZy6GjiNus59uk
5L3jXLzZA0ixU1MmpOYVne1nG/fHX2JSgA+jPrMseajUdT7EOqhL2lQ0UOX2OQd1cM8hC+Z1W5BT
v6xZLOp9fc4GueWrx0TpDd+sGOLWUV0wLC4PwOHyzUMwobfTjbI7ik1HHcv3Le313JAfzlrOIolR
GrHue30XC4QMC2kubGg2FAz0tggTEh7n3wp698mMXOJg8FvV+TA12PL3eQ7e6n5FMdgQouqinACh
RLayMig4XkFDI32VgalcAYne/A7o/gHHUfalL8+sX1hrf1qH4Sqz/XTvyc+7Lgp9LJeZh0eYGxSV
yrZ3Jhjk5kN9bNA9ezVd5Cla88aCbnGi0+dpLkeG2kIKEu+yjZVxqp6hzNFLKVQ4av9G3hLQNWDb
XF8ZJfBqhmi8hFRyFr9jw062BkZWVoPvKeOTEbbZwE3EopPSnp3RIC7A8Q1hNp2mKpRR3Z4ApQX2
gyhLfYc/E2r/ecHOkG6+YrVMGRXkOUZIzvQfqR5pGwN94gh8vALv9Jq8lKp26K1t8uyMqrQQM8cD
M+C5CAYlzExZA7EoEDJpBJbZx7KNVi82OsFWv/TQjX3bOtkGgyid3UB1zT7Wi8nqkFtdMun5R3aE
bkb9XwPw+5wvKvUi+LNVGvwoiO9fvjLHpgvCfPi5K9h6qsPwRIAEKrv3p7TuIGGlIp7y0NKogp8n
W2oAbQCHKfHcCXhse5OOx7HRUKfTqCyivXagR6u3yf/0qrnprM6hyaBcVPbngrGX65622GQCbOQk
Rs3Z6BRbLvPezObBAVQjvBEH+5n10LLABXgug4KAR78yJX195QEQLaaxa80x8GxSHBnofFBt15Gd
w6YYco2ND/vI0AcgVrzgUc7YwLZSh9ZyfBMT5j0ZEdfEAeaYlAf/2FQduqCHOfpuG1/pCoMxXvVW
ATf0xLYat1tvjR4zYsfldudiMZ9HMTNRpamT7vAJvdQxqo6BMrMoiO+LLIE3Ay+io2V1qHLLASe1
cGawWcqpRFJ6++DS4cAgetT2JgenxYHqo0LYqUAKT3c9As/1TLb0nuzMZ+AKl+MEw9bu2msmWdxq
ZZ70eUgIEC4125+C/JwbIC2G0VI85BFyLdXDkO1MRpyThIrgwKhsgQsww/y8URfaBNO/LMv79cOo
Ea8yPDyzD3UdKCjr7x1mafEOCIXjBlsmu5++2aWyviyjXBTxxRfitZ775A3eMrvf0QS/wuAZ7648
phfVvPYhwr7k/h/8Dz3jUWqsSM00crsnmpCZMOmpXLbAgH4Yo5HM19M/RLBVTDdU0QNKcZEWzbxS
C2Ng06pM0ErVmZwaUrY9Y5lLYAZtr4AWk4aO9d895u88zih3FlZOGymkzERAHVtkSLu6mFZMbG7I
49EMzCBfciSl0PBambyYPD9yL22CukkePohON8xbCKVSLrLmfI4pFwZmdPojGrReJzhfMQEaSbNT
qM+1dZ/c03WWPj3bnAz+XrwksFtXsg0TPDd4swo5SQQj0zB/SJQaKQLk5mTCVzVLJdfwdXSfGoHj
eM6DD164Ozaq2fw/fYBpqg+PNH7bjcC2BcSFl9Qq5swSDvAIhlG9pjKC4gPilIlD+kvJqg0ebVKD
RcCz51g1S3lb4Mst4OrWYLfrEW0kgOdb1ZhoHK5z5YCwpBQGT0E5BOzwUMr0Eq/FVPnQEdgeQIiM
QBAArmmeNHAxrzeKRo8SADdd4aphfyECtXg37DxaKobCpyHqAoR+uZ1w4RiD53O12bqEuqHy3sNN
GzO0C3EZiII5Exqi5fOf8yih5HNP5pD1Mc2YuHr5dpCY6WV81q4p6ckMDNAWX3fX6D+bZYol5A9D
DMmmyZ2JUvrUqoeZe3Kqs25uLCJ+FDXgAJl9pZjDVXBFTD32BQ1zyZ5+gZULgAvqSvQdZ+iVc/rW
4Guj1gyoliGKx8gPil6H0KiYRfLkDxP90xTdNdHZWZ86yRKrsVRydQnOqPZeaomMVs6Sd679Bx7s
JpikpKfp7dSaXdYX4bbaG69Ppd1+sQ5fBDq4V8TzFSrE0+sTLEaYjP534NK4pM7LP/Qty6SIJXy6
q7IIOoKRndWkZTdWTESCJisZD3T5PRWdiYtcbMD9n6925LHZejZH4N9BUgoYf/y0C/1/tVgmnlTK
2Ml1bulheaOvWMg5TG9kV3PjbgPbWyX0/MCM6Tzl11KEcpjRpdui+GQ29ttcaSQUf+YSVZHWBA8j
ZVL0Phv/ep+Spc0h+EPBz0I1iPDVt12VWFzsUUbuPjoB9gCmoGTb9EkbyuT72t80Xlq/EGcl+YBi
U6CCAJSWx4dJ1NsKo7Q01vqhmPLTIc85dXUnlrPkwH+HpNuqbx6WJuQ/gdkMasZI09snS/A2GYQB
+A0LWQPZcMVy9YEtw+kzVOBngWNJFczXYnST8rc0jbtPs4gqPC0od2k7P9l5P3+jRGvWeC27f9Zd
ZqILFh451kO3FB2awf2XNvNqm8CPjz9OkNWhocYme+BVCASuuU+2g/X9OFcdag+5ypw9F3P/Slua
6+vcU9GF0ubOpVfRe6vebKZDH8jiBIL89F2eo36ovCxeKNRYACnnGinHek8VwoyLomcnzmS755HO
0+fFaSNNyXujfiWrkd/EsoYsED8H6DC2ZW6Sx/LZ1dzqYcmencAkDoUPVaLgJcj7cjCtCbVoekAa
qa2lz5PckiMG4BGG1znRzM7tb3Eos9RQkgq1vaD0dMvNlPshpx6LzZYIswDWxbadZWAh0s/DnzHy
FCoc5N/720H/4N/B39u/60fUeXvEj5WD/+ojXyJNzfN8H3DpL/3S8vyVESPnxDskNRMEC0Z1JC0M
CC0pFG6sWXfGa0zkkZFCyEIwGKwE87am7kIS2bWSzJ7McJAG5fZFpfmtlUhplerbWfGbSqgdaRNy
38qHEU/gjYo8sV9EFRfYzavki8uWWRIAz+vU6W5BcgFhW+IO65V9cw8j5bZPShq7hoo4eWYzyPfV
2VIPzA/VVxQGrNEXoqi3DX4YtNG23ZJ4M+zAidF8/ttfM+Ie7CkQuzybMAJ0lYsQgtJwXw28Guxf
vrVdN3+NjOBzlj9PYB/Xn/XBBEyrmz54hyehO3ANpPtq1rHoZchpMfk4gjd/I2iIAKG3683NliO6
MhvW1qozhqX+Q4yoIUN/IqnKKWH3sGCJwy8r7b4DnKUeCzuQZZt0QvycSGDfj0B4yZycW2v9s8MK
P6j7jBNmyehYvKALZVEEvV3SX7bul7LUdNIlKoIJ31A34rhDmTMQsd+sc8HVgDSY49H+xKmIz01H
U4NpP01CrKtF/VUtqUUF7u7K/274PbfB0pRtJdiCwWkE4pKpEZhlP7ai5DOLtGsHcBgv7iAYDL5S
dSMFozmxkFnFREr7fHcqbO+M4Nj5mdjBvlkOWaLSO3+C634+VFJPqDkJXR5gMWnjVLA5NSpOiOSR
5yU45y8TVvBrb/YuryxbLwldAK9dR09J8wD2MGGz+ffg5LuTOk25mtLI2dexprmqslo8k+2A2LxU
fHIki8Fzs3+wOFovaaw6YqBRrGPYseVN8XyI+r/ldoLQC/PR+50jXo/7rKpg/4Vpt5cv53qrNBYR
kzu6onklcX1vSQhHMBXf4BwVNIFzM97PLG199zMEkTP8OnjdPZkSh5gLB9KfDZEuKlzQcEj0yrx3
6pr6BhgJSYv7xfOTGKG1oQmxL903fzxbM5ZAx53KyrDpYUVZfmKW7vvpVG9FfDukq11iAq4W9rOc
kEeXQbYakQISvAkH4W2zZJcjEgrD3MOUiazOIO2XKxCyC0rVPZ/qAVAbchcIxV6IijcavtgTqRcU
4+We3r6/I4o/J9YcT5RY0HR59oFsgV0LfHbmrioAkS/3tVaLUFLCRfQXuowoPY4C1+p6OkSVkAKe
GITHH9960gNnI2IrfK6VqLJWwJlTWJeOg09VTqCmaZeq6hy1EVdP/0wKbNAqG3eF8owcpwNK79Fb
Tot3vhfjQe0D5V5c0Vo/Psg0I9vF+81z+qmxGHMdT1d/8c7oqOt5FJcpcv8UgRGoizju9UDkT7v9
A8AYaDUigqp3K+kn8ztFdT9W4/y6clZaitgpJrh5Zh5/TAdkf2z5JsvPZleRkLNe68dy7O8o+kpt
i0H9uk6nD8V4w8q41RLqGc2gu1DlPJ7QUdLY+oV39oeF5nONE8uMaGt3HH9L+42/wFAKAqjfFouS
VYBmeThggvHPLdVVmr0iXDiTiJbfMrIbEhtFDwIIYOKqw6WhIR06aSBWjlwIQul/UhYytubLF4in
R1HlvX9Vsnf2j3ku8zFTFz57lcLYtc7U37Cd2ai6OadCWzT4X0qmr9IetbiW3uWPH+JeHnSChFKX
0mtb8E1e15iX3Mblt9Cc8RoVQILM6evtPQF2H328ZqczdVXqQJFn52xqS7awOcZmbwCRDDReQYXM
8VzD1DOyGvAd4AjL/kVZ4pKde4gXs+5b8INjwLfNfogaIT3B1jjVIjyxhLjHk9qDRbfgcCjM6y4A
vzMJocAMrkDunlwzi6SLFdhNAS+8I0n07DtZcWLDfldchTrc31vaQZpoQsT4WhYLNljaioIsACTc
xgQ46eQR7g7vaHJrm1kP+900B+QkbGV1N03015g2e9SJITTaUz4wOSHS+QHRyi+5I3kXQE5ByNw7
4qCXOcJOrHfTykobfr7y4i8TNO5XZ9DmL3sHeTevBovbndKRKzg5IZ7JzO8GVnmgLAYpi8qp2uFr
bWmFkrpgKWlhwrWnVZNZ/0kcqzSxIO18/kBh1fANEI6K0/ikp1URBGHPKbYI4Bz4N6DT6covycrt
FVz7beTNQxpcT7k91+g9G7s2qNVE/ICcuXWBHxw9pxWaXzoX1rW2M03Zw1PNtBGnOTFu+SQUPq7b
iYH4xsJRnOM3Z1ofU+ki4UoX3JSJsV1/cz+BxBQxEdhdazXCc+H0iQvL8Mr77W+hpWvQxchAiLsI
vFrY6fTNMM99jQhcDbRogC1HkM2t61DWhFNvHhctvQsjREus2IdH4TMZ2mxElvl0PI1ncDRgLx/4
/y3JgM+3OIVMwJ/2aO+8dYISNyfYmH5T5/x6YSbXMR1Q1kMv/wUcAd2yYhAiyGilfNV4LZdBWRB6
oCixw+W97ys6x4+V+cIZortPhsDdVNz84vzebZWjTNHZ90LYdFSixveeK5zkaj3oWWzZcZvmFx0r
b4nNWLOF06LSp3oht/XLyoVL+fHfsVSd99BuMxgmtmySBJUtYadpcncyI0kntoQ9rT3J5+L/3CYc
aGZJnYztfDgdhYLERBAMNFd0ZaSyHELvgPDlO8/XMhA6Um8mEty91ymVWcq6UqlJnxdEjHHeljpx
oUiPdcLjJ9Gkl3oXaBKMmshLM9MGegICM1PY7pcl2vBOfHv56KPsbdDP59ehkwbAslQocaPkHd7N
Zaq/u3QOqQMqsyEvdlz/2KdFijj7bnMJSf+9URfu4jT0Oo7/DohRbeQzRv/0Qe/0Obl+CNSb+ecX
PuwFBj1b4gvDMzXNmE/AcD1t45N70+IcVWSDWQeqc3hlDiXTX2xQZ22XokA38A6y52/gYY8hV38k
PEHHpWcPywyzE8DHv6gT1HuaxYsUVjBRRp8zl9SCLCWw21Ld8A/2850L7EAm1+RYiaQVALPFAkde
mVShmsQ1G8oRD4FEDss1GPGC0H+VGDzO5T7yTaZQFc1iFYZEXTtPyEtPo/rNHFwG9IIQONLVILw/
azQ4RqdzOvrs/FZYzXcK9JCxBn7MnEmfKSOacS9VTEpq3lFXe/Fg6wKFiOetOlU58IQToEoo2Q71
VCjSXsoHl2tzVgkGKDYZZTwywOoUtmpyfr37cPNmxz8b65Woqkkm3AncJQct0Nmy4pEC0XJuVxu0
YYBZXYuxbnOV07OxHxg8OJ1ljJ8Gz2QJEei+LP6zDR3+I9mU//rdpbMmlzpmlq8vCVY7lN3TiZkE
6K4Jr4sByi5H6w1OGy7sSZL/0Lm7PrhLBxfnNrGDJ+bIZ/T1kUcxibRT266zDa4MV4y0XKqfUHZ+
2BN1jYueTHxzzZk7IIHTSOpxICT/drs7vW//aaMpig1YR3C54ZLf0fPOAL9k03u7P0Xbz7hd8e+B
mUeEpuU9PEuJHAXjC78LCf/Y4Vwh0TISyhD6p1K4Yx0CyDBq0x4slPb49xERbnu+N+cgF15obIBi
lP9MeOVUb+gz01Cefw/yQBx7JAuItKTu9mz4S9jz9agzt80A6zLsNSwCg7aY7U+yzTYxtJ8DIlZS
U8KrotowYCpiW5MDDeSQuTmJNET0MjilOj68Fg1Wu21L1/FSJa5ck88ZWUng/tgmwN+hV7W+L3P8
3uvGZmdLsdhvpjLoqst1GWWuaVxu/eszYD3cKEvgU2o0Z2m9fxHGXDEfiqSO9ZY48Nn7l+NWxjVI
FWCxMmeSl4FapQYFSE+HcbVf2ZLQD3oL6RqB7eHMtEn19dd+3LSwm+bQlJDfTDMbNTF4GYYX6711
2qKwOWeDVkIumXiRweP5MgOmHphJ96hMJbhZCiuvwDRcFNtwzp4GQgnYNsKBbJwShntYhdhhps+W
CHDLX40Zxm+57YiUJ7F2uyo+H8Gz73P87I2sf1D+oj2kdG8yfNDCwM/Hyp7bfNX7KF7YOwnhVZGw
CZUu6bwDhKj93zlMnTCIxyqOxsWH+PnUrisnuBqVoXpU02fTlk8du3BqgotqktZVJaygdLoWqjwf
i8DQ/LEsDGDtcmM0foeGsmSUpEL/L2ggrKGt2aTB/5FhDttKLoSgwpfFX3ByA+JgCF90YQSva34H
sbq6Ldz7SJxjhD2BgBbW37aJMlH0QDGQZIKDxajGymKElLP6ZZ1rdF64ufJiM7+XtDPWH04yfFXP
ln6UV8+RldRI89Gfc9KxSws99opNCJSMZAw8a+TJGsTZJ4gnwp82RqIlpRguhVXpD4dE0u6Dq+HH
LgQb6aADSqEOVYsv594eouqQvU9oSUDdIg5Noq5I7v3tD6tQUO9+vLUv28rz+Crk/Tv8gH4twcL7
HxpY7vZel5vYnVsNSotue55BHEV0jweGy2A/qKKhXA4VbE5/pASjC+eYc0r31JYykBNUy5dCrHTp
n4df0g8rnHjal+D+b9Ko8vVLiB5yv+dBX1ODD7uis3IC5rZKBaFki4tyRY/gKWv8YATUM8rpgcBi
iKXMB8KSpyK1OcOPcs19k5388FkDEb5oLEN1LHxpbCe98PjB/tzwBuAC8+M/rARYpxtBCdMJro03
fGgdfjKVgryRAiLutO2aDPotb6ZaTrIetZGHZhkpSA6dKx7VuUy45/0Ka4ccMFyg5pSTIus47YAo
G9Yg/Q4kmKAvV09SaSG1uaMd3taxbGU40Z9+aC5CRqxRaLfBTDmazBdHkO5HWxf2dDcKO5tcLyR5
g92h2LyhnH+9k1nhUkNF0dDbZUdJDjtgJ6GBS8hKXUznNOn1dR+7tMjxcstHjU0F01xzBa3/f+dK
hAp7QTOOnXAwshFpwv6n0+xYGb8kc9gv0I+ezoOeUSLsos+gZFBGc2ZLt9uOWo11u2aIGhLthxgq
DgHHlkWOuu3mC4nOs3IXGsnMQnfm5/j+E90Wkw/EriKZ0iNaVggUKY2x5AGXVs/YLBytXuEOwN/j
B5af/PalaZ1AZa8ezujKUJj8d0jkcsEwzaEGIcs12bAIhUPclaZspy3JezJgH2mbuaRSXhAESpec
GfAI5cdz1UcmV4EwVa+EMwx7CUMdpm+iVdZVAiQK9WwmegwP1ytjn3zBWajCI6PKmBatpbHG+9i/
rOBNlDHatBLW3/SwuIJuABeFGuJsWUwxukpcehsug/U3YBoNTEoMuD52cO3pOILU3ZhGg5GfgBSn
rvOgYN/1AbOy3zfTEjkPPnsEkWNtdOEqOlyrNiIDSFC0O6zLuvEEoz09Cq5NxcLW/4XH0Peh8rRe
m4240y4RiT1dIXb6q/mVGjnHeZze5wGQ3kggCp7wiS22iPcHo4xbBesBkyYaDfeg8n+33zAQb3sV
AermjILv8bXBkn0GY+W9R2PQsbEnlVPag4V7TQGIFl+aKGFP7bAAcwUijrbPAyuo6pOFn/kzxSBp
MdUmH+qtI6C5HhRCescE6KRPCNAntjZ57OZjnJE8hViSE/1MiH1FDXbxML9Et9rP8OnKkEZ+Rb5T
wweQCTxLtZp4f9+hEuPfjcH9GrZvJHgHeXOgHgiiZGPBIVTvQSkyZld8BGzb/0bZzXemYtR6GG06
a5kD6EK6TWjrPPtU2aNKHE9dP20P7zolwgq0NWuswtdG2c2iNwu96eAkb8eK+T5eyYdJ4Cjm7EnZ
wltd8/7AxVDplJhPRBWTNrM6Deo5fsXL/Y4HMLp5lXApN1P1io/eWv3eXOfePW0+NFfZF73AUxNk
pE/56d74fTW3jGcJ66SnLif8/pQqwBHHQ2eTJEjwLtb+jqzz4g90kQle9HOPpLvLdSQmSPJB/gOy
LZ/JYbGEoIyFCYKDf72o3XhAHxNLCjihlVv26CObAaIWxGBXEiG2kb7xxRWFHzmx30fCDJ7QUQA/
plBk34awCCZjRTSfLbawhrZjY+2lc1wQhUhDKD4vqHE+A8bCNQgjJGZcix9xGuB6rGmrkq7YahPr
N8ElL/oVBqOTiJNXuqrvX/WcXXKmsO2JM6OqYdqTcOK+PLA3DdAvZaYuYhs3liNcqtBYEKTZJYKD
RQjLI2tv7Ji3DMpmlGSWF+8fB2t6au6NZ0U6N97wYy5/Nc5ODboCcXLbB2soWVfbm2IFoZL9CN1e
/pGjvfS4BtOPN/XE6g9dS0Bj250JT/eo90z9jZrH5T4nwtcLAndE9g4WRWtVz1B4L6/QMW9WVGjx
KGcQc15Y61Hyv/lCi3hoeRnd50e3imoLN+p4EyTTUksN97OyFIg+jGqRPw9fkwP8+R2UJck2ei6v
omjU+c3EveCN39h2MH596y1ZZ/rcFIIqOFw0qbC4pV+ilJc6wnbd0Vgu2uW6jP/RAU21Pxgf8R8K
77sfBEejM41NZqN4PXyaq6DIHoBDrHQsm5Y0yDQ5LGC8ZcX0cbKcwKwy+9n++Oejo8dqoyvUV+1X
xnSJAK3GraZItyz4jOCU3XVKATskGFBdzWj6H1w2gCizOkJ9QMfcPvHzoO7SsKeZAUZ4G9VJFl4a
Dfh0+p7sPISu1Xjs/G1LHVr8R70JNZHcHIJLcMA5s0Yh2nRK2q7Gbe5IhAet8Faw5R/nR3BAUxVU
W10/T0f6ms2vspr7s3GPHlNc/id7AfqcbdlRNloCGylVHwyzheeISc/eolWwGU5jpRDdIShI5rpP
v5TE0dwGTzkSJKlDFLYi17Ez8iOVsduV+LO9LmJoXI4fTLfy2mABIhRcXyapC+Lqmfz5vOoB4zF3
cUoakRN8TsGRN0N9GE1uEoIr4STYRn56hc88hWZPCdzC+rYFEjmkoD7MB9o61yEDJzi7nxewfdgM
SJnbz6DEZH9zvAX3IIaPNhJfPTx/suh8A76ta6Yu931T/MusNJ1GtQdblg6fwPXGZDOvtCikseoy
5IQrIH2vOOx6p5AfisKd5R5+b1VJl4ccDj58jl3hKdYNS+/LFaDXs0F2ZR35UhlxX851ocECE45w
Ker0K6YCsWVq1GozjNAMS8G9jKF6GRUy9R6ptHqM4g+X9XJosXhKzFtTqy6gL4tuj0MAXCv5yrmj
vfG0ymvcMG6xj/Qiv9CTH6KhkSuuAUDUzCRDbxHYmQgy0ij8KN3n2WRdk/sYuzaMAZEH3WabACTi
oqWzjRdvZpLEQow88IznqLlnRZrgaslKjtl1TWi3uM/2t4UKNE44ByqoODjXIk18V9/HlZLv/BIE
W4lzYcJw0s1EXZoOhQ38GP+ECPbmPwJT8/lXI5AFWuG0Mth5e7MCTXkFFnc8oTPSWADsLYQjJcEY
Oa4fRK4OzpXrwMRvERUBqzxdkMxWIj69ybW4RbF3jfJNFeHXlz27K6yAuv9cfY2VW99JNZkqR4ys
ZXb2m5SuqyYyPjDIkSbzwENzONJwE2gPD8GXFRA28Vcc+yR/spAsDlRZlXa/b0ZqkaGumE9sldQ2
xtRk3PU+V8vg7Mx+T7iYi5bST4FdatlrcxNwQxSgIozidjSHrIMKjuMwkXRKlIda79zq+N/+Mg/P
hOuBZZHojIVbyrNrSi6MN9/5EXXYL6+HuEi+JwJD4XQTVPmpsUuXhE0nIwjO1Uptr8n9XolPnGn9
KKi/jy7UfYVAnHPKu81NQy8gFlQC1UM4Wraecgzm4DXLu3Ulx26aDx6WNuEcxIynYN21Rp7ezgw1
5RX9E30o52pNrb3IhwXI9pWJ/kEH1D/7st4BR7OtNCLTqJ9p2Azw0lBmkOuiUfBEH64/rIwwwTvv
PmKcF5CEuyzz4cIkSxs2DPqcSbH5P9IU5eVGBrsNDmS8t+yRlWzFelywePxlCub3FdrMyVwkvcVX
kJug+SnRHM9SAlGIKBu+rqGhnMMTE9CGphgzE/17wedBF0AZwyHK8eg/Kphn+2v4Yd5FpI6+qCek
Ct3qTb/cvmX1ZssreoUQf5gCPA8ee5B6eRfBM08CDVURcr2SpeXrC/GQyNB9Ift+qyd2i/La4GqA
w++65mIM3AKkZYS1qnmr/3sSfkQzNWbhI2wkrfaXkqCW6wrSGKEQbrAsSFy1B+HPSNuKCwQ89QxS
SUc4NONixoxrSsUIAiUdplvcnvSB+je3BHNfn9xxQAvvTOICpkYynOwHYbFT8UIFCmNCf2OPSqVa
FplRDi9jit529rksM/k3m+zewN2bRrqIHy/ZV5Tt66H69RvVzGPYbsDr79J4zINjnf/JW137qby7
Z63RyUyo4O8avkHBBI8Mkn2q8RqWxQ5uy9oqi8SxjaPEsQxnLkkr0myQZm2dAPSwHJd4ThOhAgOU
DF52/Zr7dtgj9ym4PsaprSXrh5S2a1AQ8g7v14HoYxlIXVF/P6mAmMTWwJ/zhWlhm2dHPm8thEo+
kPB/TxEoLtONVu/1MkzXWB5Bj6qxq3kaG32Qx8xYB7LCCm+ocMgy/7eIHhS3XXIhrkingkC97bZR
zmBGSDEC9BjtCyVUVixMYvRh0A5alvr7Y0m6Jy78oqIXq+c8YhxyCv5/EvC/z5UuxxphzkBnSRXS
EQC3dJZxQtp1XFCNC3kDBJvNXj7dG9A2Y+JFCcCrzBaJIHYzbQa/e1KTHqMVQhQnBL+hHkNeCl5H
dOf2BzG8ZKiU2lZGI4F5zG2unlPlpHJkIrGNf+Y/2EoVHlB4/+oblGSone37bfGv4pXE9zetV/8e
pD05myZ8N3d5VbYrbLV2RhbvWxXhWwQEFCSfcFKWRP2mcqXkA7xBaBIALfe6cTzvO6QGNcD7r4mj
8bq8ro07DQOMyARthuCB+um/JFVhCZNoR/73ephXAN40nyYy1tadRGiUabt05KIxF2BPwsAeLspY
0vuCxT9bmoH0+tX7ROF232MvxjZPAVcNBhfIWjaxpOVU2tc4oiAEEXulkpV6DMA06mZaLJzFvQIW
CuN2YtnkdtFJJebGoAkDcNbIBenkh/bMrwJYT2jmRuHf3xCBycfalL01nqezsdD/UBm09QhsKHen
wE5qChd9AXaL3XF3pwHVtZBzHFElmCBNpD+72eM4GCi/Rw7uwccn+LY0KhR2EIrm3o+X6e8NEfIB
2bPHRcUfFbnsqrooOm8U5w/McBCwJXAxF67zY0TE+d+isPQdtYo6nforS/RuIk+aCSpRwbn/oUY4
KSzm/XjkKG9NgNMIODkPdoWpCfyDADUv0cAs2qEY5Ze3AeBx48bep9aNEJI2rs2A6R230QHxgcvV
Ru6jaMt+C/sB9/TmzI8ygazZsYiO6uyWsC9Kx1BM7guKa5pi0jht2Dpc9zPVdxty5jDpHtMV5aQ+
V4Fgfk0u8wyHxXB+u5wrlIxp/cRWCVnos05tn4Je7NLaZFgk0q0Gg1+dE12eypIfTzIyh+gh80Iy
XzC+gd7mQeumvK30pjaEJeIAmQTyCPaORsnoIJMHM6/7XwuQZTc1/hkruXh2n8RVnxPL+dXu9QKN
rW+Oc9Mgbw2QFH32wjhxX+5WUf1J7XkHUPCNHXM2BJTx9dEJHAmxWbCZbnL/hGx9MQHBeqg1itym
cDn2JtK6fsfPgu0/jeBAWgoy6Dz8wPx3aXuvMJLmkHtWjI3mIZlWuuI97LEGMFbqJmWsthMSc9u1
bC3WX7cZN2at5eWSYrogaftaCV3EtDhpCI5jxuf565dIzDfwPG7zJ4suNWFWhVq/Gd1pxARkM6QI
5P9iC2BSFIzJIGGPIzW7D6Cqs38ppol0POD9Sob4Z/QRIaAB1GyS/pinJE6ul/md9fNvSlJE28CG
GXUvrwZ1i7ZgAq7UXOYw3IlLRfQ1javlAF5KosYGNk+kBh4UjSGSOR03ThqhWLcKEyvhKz8WnLvr
bPS+XCj8duyJAK0TTApf+4TX2jci6bV3SSOPyC3Y3EpnSgKDz2t3FSX744mhxqNDZray2WKNJmUe
bAmKL6J+uMlRcY8hGQRmuNXRH9opcYXA+Tsdo5borZ5D8tPfwLx2Qjkk7rk0oCzTi+AP+mOivAYA
2debnKkoYlGYrXDuxF4XSnpXFAnWOEEKefp1KZi5GZLkOjCdLtP4/c55VwF7pH61cm0mO2ppI7XS
saVD0VLJwael5EBj5u40ZQF/mfslzKl9taYfEv5HJ9F3qdX7qP1P3+9sESHfh+np1wOAu1SglRAA
eJ8yY6BDwhnVdVGkMBP5WG1N8x2VkmemUtTa1Jkmteb3LSrqEOiaPAToKpbS5ch6aCbaaE0RTiiE
JucQeosRS3bGxPW+HKHZs/BoJ2yIXLuQhHCs0rFlNQCGmFFlBNGfNo98+ZQY6Sf7lVwSFrcIshyv
y26pm8VEmkXj4BsMJ+Vg+fW8JogQlVrGtv2/meTmeJQhE9g/Fch7ljGbQCFJklIo/88I0YCJQsDM
1fdGdpa72+cfbWWYEwiIJ+YSh6MgQRfs2ItnnebRelNMH4sbMeUIS6rJYHIhUiDbEMcjWyVvTvgU
zE3Esv6BLXiXjO/xp2t/7rFkavY6ZFHYAINVV4ls/X7SIeWebUVx9yAwTWV19iUKADeIoTIgR2IW
IgIrSb/wa7JVexTnbih+5AVmvIyILhdeAE+nxTk7VFXBuj2VhUS0Lu+Zc7Y2FnfKvwWlxpKcjJWv
FWUKUCaRBsYtWt90r9aVX1WN57gF9blEHpzKi0xxIb98rZRWUljOUX/NO1aoMiU102iDteKUgC4o
uwlqNyq1zgCWYKWBtO/lkPd7EB90c/1MVVRvY0ruRj2OD087/HrgV55wUIhByz5wQA18QeuDyWi7
1ZYBn6o5uQtLNGjkwX3vUc+jnGla7hjlr1qXD7IqZgK7UhvI06nM3fMNGIN1A2zs6jjAuvEURMCr
/Rl+yC37KXJtuPpJ/OXRXpc8febO0rcDD6aNWjps88N5N4oYazAwQRuL+zIZ+ERRgV1sL4Lk976n
OW/2A375qli1L3CqCs01EBZlO5ITD/w8mWGvtiIQVz/XrDBL7rFR8WSgy17SbcmDChWjLePKW55e
sApowHQKeZKM/IoOF7m/qjATT3Pym1Hr63M6eQqwTF2BFAAquO5aS7vOojapswMabEKWD0owmJGr
n0Jwk2ndC+vGX4pTC0yIFp586kdHTm3DVPAMgOuXUNzMW3zSRpnLGFhRtXTeX2mapq9PnoR98hF1
uMxmVLgfXFV34SXzW7nPfpv41Oa+l6RIiNkAQ07Hw+mPXxUcc4PPiUj7uAU1ehdDCNeWM4arjtuc
DDSOvc+HGa55lmAt8zRx6h8nwN1LWLpYyJttC3PbQO+rIme/FwxoacNB84cs6AfVnv8Zm9pT2R7V
ZDwvJpOI3/mRodfw0+4zC0hFXkzoozPtmIDj24wyQIXz8E2BH902g/fTACfhwiyBgeoZI8Y3FTUO
hke2jVqL88cDogWB8+Mjf2yhuneQYa7nvG3UeqOcFgin83HUzBICU9Ov93YDGYEXEd4WknNNrGft
d8do3WP/NI956CFtFwdZyBjZegqLu9Jlu1xeD8hsXJh/VGF0p/TPNzFNDda0YxFPYEYhynoaNPaw
wbW18nSjf8k5PHJrVkbwUg3/6TSXvHB09Z3U+RdS2XcUlF2tK+KUdvaiFc+iMF1oeUdgNtd0tDhj
XQfKBAUko272ruOgiPPNEXUf97E7Mb5aawmF7CyD41KDudQmdiMb6K2akaIsVZ20Ztjtw3AW29vo
tobt9ilcHBS+cNHEuiH+bo6x/BmKeV60L4qS+SdKOhu59NU7NxlZygcuj8RB/ytjOvea9al6Js2J
SkvHUwqyBPDZ28MtRw5jxYOiN46R05yPxSLuwy3Oz0O9OEIsbEcgbG7yYWXlKTFKI/p7UBd3cdYj
9NY8NhSxGcrwAVOe7cXLanqrWisfac1392Td4qUIskpDtbLqV7kclkRdwcP3ubWxzyJ1lJ3zmYVx
jCOrRGd9JddK8KOV8GxrD8a6hX2GNFvAUDUiklCWobEzEo4R14gR/oiV7HKpFVHizenGzjUVOKJM
3xho/fAEcmXVzjM3qxUTvea5KsHACF8SUAdtA57FC4h7pTm0AxRvQb4f00JaPewBUWkmULzmPUTe
qeSWd+I3/h8EZ1cLIAC679EHuGcP9yUWvhCBYt8tvQZ1wCIeq8o7lpakD9QhRKm0PN5xHSJRnodC
t59ulDMS0VqlO3P3+3y2SfUCy085U9aDRek9dhOTne+iy6VqILx5IBNnUF8loXHBgGYOJAqU/Yql
cvCYma4xqGH5JYw1yuOTpaLv94qFnJCZNaSBNqGi6hHLy6yNKB+hkVlDpaTYRvUuHnGyX3Q5eR4k
FftkCD9GVojJFufwMlF1bKSDcx/YvPPvZi3znH6ghhC2+pllxm2ON7scPxu+vlVMEvT9AKJxXwmW
dZWE43BF4Nkt1yj9z8ZC2pmzRZxPiu/P1CmRI68i3EPMvjBNSdyJqRkcRo4TgWEOJfZJkhLA/Axk
r13tytAi1RIVr+KmQoacRbeG/iN22kCpQm7X2/LdT4I8wt0Ry8saTnwcOB9lPVp/zVNn2pSqi+gm
tqV1Kssae3HXEfXH1AG1OUYVa5dbJs4xUhh9pPCsy+5DTWNEVpvbFhMj6728bKGEmWvmmLmGH9De
bW08Njzy2Our4fc9WWVjU7zRz7LBrV7sOOJOU6ZHrKLSvHEUFdaQs1GfWS+Mvi2Xiqtt1RRL+6FY
8mawai+k8d70FFEwnA0RrNFLi3ZKT563Tr7l134nG0VdN6XvfI5HYvluq0JBPmdJ/bGOt9MAcEMC
hnmTpeqsbBsWCCFlXjhsAC9yJuCI0NxzaClN6G4br4U3eiKo+vTpF6FJUuHFOLuEtBf53NfkqyQS
qRqPorJwrYpAfkNpXUzOlUEXcYfkkXNzDJQZY5Mu3Ice/uVLLA5WAxKr/pmZ3fDh7RsguODILeCr
qF6z3J1NS4QGClGIjE+1xB+rr7NLgWkmDq36MJikAQ6nA/9MiWLuKMK1g2eQm4L1z/R2VQkAISL9
ERqASHS1OHptJnAemgm1WCRYR9ZBSwjks3waUBp+gVqXNBG9/DZ0l1IDF1xRYQEElKePDFp1tGlu
pQeYjNHCFISwsY6kbD6HnV21HCaa6TDlC6oBLkfCztwG19asaCQqSiz+SY5MHQ3sIZZH8urwhO/k
rF8GGbkFG9+/w5NBJ/+fmTRN2GhdKfAzcA+N/bIwCR0cx728ukJEXc7ejao4stLZSWD77mpLAG67
KMSzo0adN0DTFJc6GFTrMFDTMYbHKI1+PdWkzFN+16E3Nd8853El6xxEK7kpRSwjtjJdUIObVA/+
WNNZF3wQmLxya/3Fr+NU9WNSOv4zT5vr8oTV8XxbO4tmgInHrDLwGIrmtPO7K+bU/mKkOqae09sd
qqyysID7UBtRIepr0chK9BzxN45l49jPXzxujhy5eBLnFNBcBr1orUGYS3PPAFDHU9QcfmVraXc1
7NXpgOJPVk//TW4/3t1tPGb3gbL1nUanX7e4eairCov8GBIhxODCd8aB+bxBYqhF7800h2LPSC4k
lft+RmicZFaFzD3rQelGzUlKalZwAJ7aiOx+/mZPMCOj4X1sBl4fVQYMSLjZrgDdDN9p2+4qQ2H0
N9rcPsPUa56r5nwHzxAGT1lZkCJoX5THKFKTSywHs+a9mSj3s1THGUg2G5Cw1puazLGrC8e8NSnh
PS7kE92Qjmv3ujeMXq0u/lt+SRx4iJjHmq3JgT3iJAy+N0b7jru7cg6Q+KNJ4XRjAGVqHdy4fnSm
5Coq3If9Z7c+DD3vyr91Ymm/hW9arXKVTf+1kOBIISEHTzsv38eFQfOwv2QMgUXlzbEB3A6O24zZ
a1FJaBrERXdtXGTdhjf2BN/RY45w2wnkEyUqxOe6if42KsVaPQ204tBvc3yaAwRZ7UB37/8uNPf4
ZsT9vUZX+0W4ukpBmKm9McW+y6JTst90EpVRSQWvUxerLJHB/v9PJ5R8UAvDKceEWmC6ili0AWAX
DWgrCuplctHNT/ScSicnGooW02VE+QMpWtCTSRb49v35y/tnkvt5/woxgMa9L4bOECYPJ/9bgCKp
RWGaGPZ3PRMbHyYrVcnODGfGoy/4k3xPM2M3k5jgoa43I6mtgnVF6hYteAKNdlXz8IRDSDiTgjvj
7es03tfSuiCM4O/fGU46sDticGO1nZtqmaj5mwqlyC1vTRJY6KH1EcwZUxcOxRnUZmcxOgL3qFbD
i/B5BDtc1dlDoNQ8m3Emo0Vp3SXLgWA5B4lthll4zIyEqxO/O6i3a1Bkl5wKkgF/m982RhUQvVsz
wfnQ8WWGFf+u4o0GBEyEG+BW3+dmygrMwIXM/XfdDEU/C/f41Y5VxKTbhcRfMg8gWe3/aoyQHRjj
jU+UISmlLAyzDk4ElvXIY+3QJ8azb7A+rAkljgHcs0Hj+InY1Ynos3oZBr9ayUPDZt87SLk67WYt
Zafw+NATqd/btA6hA4gdjeOd+joHTD6aegzZ1oIg7M0/zA/mNm/ucyH0X5kgdPXRxAgjH39TYT42
wjoW9jsll+fkj9+drxD7qOv4YsSei7cZx0o0qXf+QN7pAG9UsioUcogWzWP+nNt623XuIonBCnXI
QuYzp52KnllPEVXd3tsJNg9ZyGeCLX5xYqIIysy10JizyT/Kf5ne+PzO4NzhVvS94o6m01HwNqYY
FuSqAVygbbUWCnJIelnOgqN41Xr5oyPgCPPEb2GP/tu0aTkOAi0wSS3eEyYq0BnpKrBkPfGG6EXK
IPfW4UYHgJ06usav3IdwPidAIkIyR4p5hCst4Iik7UHzeiSvxLCNZhnzwKaEQhdHni0Clste6TGp
5aWSH47wdpGlH9MFiXzhpH8To7YeeP2VhK+9UGB2PwKZ8DZ2VxD0lNA99Ck+YDCVySCbvlZGSteA
vgUgAquomtRBZ111iK6hVEh7zSyCyqPtEYzaFlH1c/IwG8jXFObTzAQV48opOlfpidKoqyu/beAF
/0FF4AO5E+QKn0cbZwVK8iR8lF0aldBmyUi20CZNkeil7bKC0KPPG3RhyvhDBwgaL3/QlCwaC4Xb
7gxqwcqCpk5RMBPFvp+hFnsB+HyGkYR8n+0rRKUi9afStJ5NrfBGUuoQGuToqI+fMO43WCM9EIBO
cpy/hBVFO0qU9ZIHSoA+cSlnYHJbOLKd1d7IJ5RVqvuukQsOYrqFryH+GEu0wNXsUcdoux3PDewL
blfVDPTpF9g241GXG6gHgsV2a52GwupainkemwRnx5QVsxprhEPzG4cYdGmGs5LUeuBkbmXxoQLW
sneB2ZN3DVX5/6sf+GW81S12DcBXeIvORXVCkNQwKU8oIe7JgFeQfR92g8rkYVk8vXyh+fHO4RFa
M7D2QXUw9Elz0nArAvnN91p+8fpyx0UqwvnxhdSUO82CtBVgQz/v/OUsp5be3us6bBpmNF51jYuW
3O9EcS+Y1iI8btFkdsOQLBt/DfNTTQJo/PIu8yr68sqSTV5jT4E3Q3JeHf2mri30in0lGtHbNM9p
jriaWOTHEiSRseYWdwyHZvGHccFf52gY8praeYiNsCzb8j7sQUkHvYPCRlwRYls/Zzsv5twElRy3
D1jz9D1W7cHY1dPEvTpbSHbsGAaNBRnQ2WgGRfCSAoReKU+GiCwf3quVxNPekD8UYlb4LqgSK1lK
9VV6NEMivhmD69VcBO8YRVw2oKVj5Kpt/pEHUFhyMZ80I0onOgGyr8sWr3FscZg6AaKpbGrR7kzY
yggUIsowg0SLIGo0lyT0awYiAtfdqh0ebOPNT0331bFvmQDdYaz0cVgx+4q9ewAtW1Jc0XN7UVvi
qYjPNt3xwdMfqY+IZJ/TOKkqBfLaSisCFWd4uoUT2wflv3gvpcuB+Gc0mtM2SAIUtJqto17FafnC
UWv98mSyQLzGgWwJi6Ju6+q6Nc7qr9VsTrBOlbhDH7gwlmUzTVfKhgNRblxwFGSrSaBEh8DuIssY
M7GlJV35AC5VRYqxMxW7M405CCbpNcVkgjI8jWVpSHZLCXue1jcMdB783kf6SECGJuyBJpGAWOZa
FiObHRkkwMKo6PXCRMXLwLV/3RiFhV9NAVKuDspMw9AI8mw8eEv8hNfRrtKUD4Hte1Cx3RjjvZX3
51ABveAc+roVv6sWOhBdyZ6WW5ec7RptPU17rpjwLsdlsC9bXMY4rQXvhLQwKXofNA9W7O54ztZ/
KisXS7mO8aor9BVzXXBWGGSYlrm2Gb9IW+bpqUOK+ktIsIDzghZaFitbNM2DFXYlMZP8+9RVq0Bl
rs4su8NfhQ9LMjCkbL8dEezPatq/aPhkynLQrxM+umFjo/PgXKqEau6ZeczTHO6Rp3GiPYCqgjgP
LmJqPNnnkefsrD8Ke8pdXUkSLeevO7yln6ENCmVk62Rzdu2JlAZ6f/WuBT1WHKWdLazz1Oyn5wAh
pf7Xt7gN7nvDFCqeT1qUImuK3WI0l7U2b/joM1lcq5oUEdm4aliSdG7ouepgv7qeiCR2Ciuhqn8x
eYaoZWSVVGTkR+XRKNwiXfF/pAwoD1LHds+7FQ8/8CN0kTHfvEYrBoIlpa6chAeGOqg7Vl/cyKYm
RgRafl94IZqpzjU4WSXDfpycygZEN16Hw2Jtb1iZtiTHSX9SYorBGVy7Zr91gbuli9/F3AOqTdBb
sjromUq+6wxu7CyJHYY4/B1FtsTiNnaBL4QcCsIsgoD7vKUfQJpfIm74D4P524OWg39aNNKBrkOo
5uHtRVPRKa5zc/FjGVIx0NQni7cgMP9eU5Ux5X1K36XwFbpPjn8++QwTRnEEPxq2LNrtRARGCe6C
abUh6s2hOCibrAXeYoZ+khWmd0gRdTO5iv52PRW4GL3lUiK4HB3qG++xHVwDRE+VDG+GfcezvHYT
HJZANrH+XAcLRffAJElUdRp6VSH8Mxl7CAyF7A8YI0ZGBfsT7RfFGWpfmD7qcKQjM3zqYztzXjht
12vL93zUf1QvPgKj3JUF7VKeSjx7YBrSOWG4Wqx44KSmf+r/znUImPeLduNPTFouztHJ5NU8yZOw
AdGjX0+5+UToZn+1b68E7/bBlzZDt7XbvHU4wilMaDSLK6qS+tT0FpsZ1O25ANIZMDFPI7fOGPNE
4WZVWQ7inm6hh06xz65wEtX8u+kFudayxAWQdV3bVWmFcrLwhEFFxS25FRqRi8GRovIcEvzu5eF8
rRtrjalcc4OEfjXfWvv4I0ihftwMX2rKB1jYNnbVUjrgcNWSCFyhAOv9inmRArFFOJV1SkzatZyZ
sQLhndOrxDRHnBsrF7lDkLh6l7RbQWIlh32Ly6zLzaog6jozhbUnQZ9t6Xqc36c+iONb3IDNJHSD
oj3ioADxPXCE4NCipZsQhLEC1obOmBMpsW44crKQBN4WRIrDxow/H6dtsB9Fy3fJcV7wSM9d/rrs
wUu9Zi8sNaqrETUKeEJMwdYIoWgvryD4e26ueitSwT25k1EaOnckOvDJKg89mfd0vrQRaY1J/6G7
yojztuZnp7v3yooDBcMuCW02X/z2s83x7qQpfvsgcgxNSfWxeCim4tgdAcEWLmGR2af55umYGhrl
rBu0XGClFfEu0MJtSt/+WCumUgjORRwhPCuFQynyMA638t5wG0euezDh+4CLcG/U4F1shYUHBE8j
XzByOfujYcxiEiaUdivmKIMzeatj8Q6GvC13sjksHQK90LHIY2RsTVw/ePB35Buv4DrUuEk2bMhv
pQwM/GoMGkTxKwVWuvd0IVE8JPWaaB/+RktTWhFe+MJwUnq1L2bx5zT1ZxEb1TGBI1wnRsGNtmt4
r3hSLwGMQruwNPiS9il94KAWZQjyyu61co38nv7L/lVABzH3Fxt3uYJ3tpOpePuN0utWcUZXSRY/
7quFr8N3GjC+QQ8gKP//v4abe4hs3sUpxDboCSr2BfJM1ZfrZizifyb13T+2YhMHuI3ouJaIW7XK
uwQ21L9QEYvrhF6qe1f30rYnDt22t0mEjiOt7zliGLDXOnD5sAL2sSgqmGnSZXNVcM4hhIsxzleC
32KmIIm0TWHiSrY77mA8lNcfUo4Iz5pAKbgJwUDEFALpXjz+ABfaodC6gNmqHWIgfaewzBpS0Q01
i3dVIGSZTQd4gc7D2/ihj07cZGOrUxmtKnz4eMRNSHxfICdznfNRnINEwCEOLm8llFlr+kW00oKV
Z2R6A1o19fGj0fwUP5CQP2Z8bG1jUU+w8IRa2ZSYpyWddFl5IiXyUouAVUnu5q7YhI6/gp641i1g
sly/Q2uFnCsazLi9hxHL3JmOLKofVYRQWKV8fYeys+h7X6Vr8z/ji799U9Y8JftnZobbCzq2lC0U
XZ/QorWaA+Ah5xBRqELpJxUeNc2mRWW3iukwU1PD7UQwykDlQLkz+QpZDuz1ZfYkvJDJi1XnhqTx
RPMR/AeSt40reaQ4/FBwU9ciRfqS67K4bxa9eWfJXAF4MAo6n8sXE1BbuN5rTm3qOZxmwAoYt3YW
gIJN5fKnG1mAQWs+O5WYSKoHv1/RJW4jtgRnQA946a7qJJPPzKg+DK5gS7SDFupadUlij8TkYkOx
0za0HG+lOrgJ0DAJXBI5xOmrDcj4GgB9iGnm1VZfiUISPVfd7JnXrCQO7DtwnDr02RXZnMALwqjx
MnIyPYL7qciTW1cWBN4sIT5Eu0JxsTz6Xldk9Xrx1VbcCXEK5flbL4iWzh1pQ7VCwjjwtkY61muL
NBWc9lfLCdyqTYP6cuJp3l1BWxCS6xbfZnqXlMciXhJ7d7VLH5MALcXXqJcnDac3Duxhsz0H75M2
Kg3fqAbBiYKZWlyb5VXsCxcGRLQY4JzUPVBOOdAbV60w/wtM7/dyv9ZLVtS9tIhUvOg69SnaD2rL
Pf2CrcmEfEFV02SdXaN+VN8tIh2YbSShqC4MeafLwZD8tE+Ycgsex7yb9Ypc3UPXqLoXYK4cZt5T
q/HQnJAzdnQXWAwnDKMojJXmnFdibUVoRJaWxucVfrkV7MoFSKxnezKf9/iWFvoejmftu8KJzeeq
J3AT+wvrNtTdT8UeeuXEa+M7HBQOt767Nk/lSAE5sll88F5ebLwmdxY9Dy5MzC7OBGHLsxsm5VIM
DST6pMVFESQL4DII/NbKBbN5SrlOCdfB8UXicXWkdBtnXt3a1tm3OTpaSbQFJGbOmmCu3rz+sSeE
tJx76ilRvgkeIHjmAquqoL5r7A7fTWh1hdoHCye4Xm5OFjxTNh7ruIK/i/AoYoRIcs3hGJAnMoYx
X3ap/SGoUOqYi+POEUgsHBWpuZliStebN7V6nDQpvxxneLKHxlLoqUeQ5uG2oIXdhcruV4ioo6Fe
48iiYDYnh/JmzqZM7w+edkfAY9JxNWKuRVT5oUOnhblilr39Ol42DtErjZ+lBl64xrghlQc1waxM
mvJNUN8aCf6KVR+R2dg9GiiWPhN/zhC/d3swtiQSugRMl+SqE8bBcdGRLhoZm/tiAWJiCjSuC/0K
XSRBqcwt74mSnZnHcU0Z5lILhWm2qrTsH+mP8Oecihhc5866TP5ZN+eLemlVkilYu7kElJ/4D0fq
m+WjcFyaiIssjOzsVJTOC6e9wJxdE4ZlNrFFmMSbBA+UaIgF08q8PSYqitryChTUc/IEHZ8Rvwd6
sqeFWDOHH0i9mvNZRPrU8MlxwYWklFlQxRnvAkbGW9wePaZTSSCB2i0UgCT/HVwQtgr2GBnoxnL+
s0pxvb00vpCxm9IZouGpqos9SqTvSYiArzZ5ofmffK/ybJNWk8Zytki2g7GkIRaXTqPHsx0MQVf9
M/tH3tHoSNjlXNE1mWayWIOHD1is5YTPbpff1krm3ah5cHweEm1v1bTKt38SzqZMRGCYxaEK1Gd+
N7UsHszrZ/WDtomQ27s3zwEqwaO4TSzEUwK6siBtMuHlf9SWnHL9JOdhwrqwm8DtTR1oH7/K+qNB
xI2J0hFd89I7TKzhgDcNSgFRbdY3vttW72ey61rhUaSdDbq+o9cKvFn9BscEFYyJUj0maXjc1FGK
I3yw7N2+xFs9w9wyxeZzoPLtHyKMGMBqjbJyBQIdN2MJfuUo737pIyNsk/GM/zBoWkdZUzRpsK97
lFHzrBbxRKg8XD87tYwD9/WXg7vWKhrAjnoTJ5A1RTC3PK4kQOMaBwvCfDN7R3NqpRMs5Y9S//5h
vUTXbZIZkGPql/fiQLsv6PybQ2D/f7+0my9+y8CXIobA6qCyz8KGZOHG2EgAyEccSlEmh6SgNseH
iQZy70o4DHoJy1ruqmJS6WiyExyJ3USq0gSM7MI61mDaXAgo1OphFRBlv1xS0A/2S1jRMLyuJULQ
50cawqRX1OsvnDl4QWnVFX/E4A7ZHbI3mZmL4+QhDMtbwJslkATnr4hyUokHeSM1o/4GoV5XMgf8
JhsSb5gkrARFg2zDcZrh2Ri1x9w7YORG1xn3u6D37gBN4UhuOyxeU6h2Oo/nwsN01Ea2Rbq/V7//
MUul6tp57UCd6kVYmU3+G1c5LUeh/qCHcftZPGNzGHo/lS1SOrN31IPZHBtiKNo/h2MS324KUhmq
pWI23B0vrisihTnU207d8J5Aa4eoaaaQQJZOHoy0r04iCrE3uQTT4T/boSe0Hq716dIWaqxMnhBi
srqg6EqD0qb9EKUDuc7dxwrgtP62YJ9n/5C1YgkBdznqYuP6A33kXCs9jJyNV028e5FyRXqixByh
duUstQufr4DidyKLR/lQcydMxpos5raFO9eLu8VfWMZPKgzXUBtOU4j0wpg3P516UGnDeD6LkfFk
gpwgMYtr+FwtAy/GrGJ8l4uhc2eVTAvt7EQFgMRWNn/ILd47IEZKphl8rvnpYUGRC51xELmNCZui
qhfEY/cyF4/WjeMDTqDkTdDVyMh2O/1Wjav0wZhA8CmFJwLtdtRZwgxTNEoCQhYJlGoKZPh1MIbq
KRaCwYV/BXfETAERSDx60FT9Fs8znKcNvoZc96TcUk3zDh577Aj3Kcv7LO7PebP6X6obDhs3vb1C
/eGbCr6fOIheuIMJlKbVfsyt/K00wvFVI0h/s7FNeQYT5uezF72fhpG2mwJJlF86ifpxLd5C1ejN
VFd9jq083SxW4dOR/D6cjcH1B/VQMQEB21xn1yJwdbC5irlpwxQzigedGlUquLwmhrPQsZiaFdqg
EUteDhS3MOqUU0IXLpZoc30WLAkcdVGkY3p4x/nq5urvt710aeNizhd2aU14qoNlZEnVly9PreDG
0AnPpp1W0Mqf6m8jbrSmU7s1wbglQLfXUUQwBeO64VGCQ0VtDVfBhxGhgy1r/WW/ECMPsrdDaaxV
uA2/KEEhJ9tUpHOm0eF3kQZHF1xp7IK5FlpwIBONKzRBCg8P1BHbu02wLfOj/CQCag7MS+Eg9uY2
lylMvi1b5go6IC42a8pR6aUwZijpFR/GEC/FsjBjbUwYPf0t4wJmrW95ZFXYWyvP2E/sGi6xwOrC
ADEYJcs4+yblBw6qcE1h3TJSWO20ahIAqOcjxMZMGKzCfhCNyB4wFsm9x3nfMAIROzTlyQX+s1LV
FSy/YSEF5kZwWWr+Te3SUr2uvg6x11hSUi7VWSMK9oOgPT0SVIezm4He0owbx3Hn/4UM54EPGzT8
HBlSwW7lkJpYuTm49wab16FGXzrEFztDZ4pjM3faD5fnKFkQ30MU3rC9B8aMNIc8+u+yEdpA6K9w
Gv9iyVLfTxLri1jGu/M73l9oJRLOZd+7wYJGgCEvdldfwhslmGEcqSxs8RlnJ7JPrpSHfRlY0MhG
pMFxhGy4y2FRDg2zHfV5V+bviH4IzHSvOJiTYLs6ZB8jdiQLBTuLpD5/BA1XM3rkB9kMHXHdVUYQ
PvpCsLwndWVirarZTuic4MQMY3qIYoHu8ZJF/SGXhb0BT4xfhY2E1V3841GzxZVc5XUwopGzFMTd
z/CG+HPQvZftPyWY6Cou3enhzoPxMEWxZe9KLQSI5mczbrGCQ4UjkivaAdl236kBjzDSK85hwDCv
qj3cmUTD7y5HQn+AqcXqXT3iIY+NMpc5hcuyOEmr+aI7Ik4gGvSRP04Nt8j2cH/+0tWcv67K2YMN
rafyvrUeXD0CMvo8y/9Ssgpdtn+mvGfIW2vUusYfYjqJI2vlD4zPpwWFp15T9XBtJxioz5HXJMuh
nniNN/Cwq75/qvJAUbEYWT9IbsZLzB4KW8bJTEOhKO1Cq/Gyf621WdYFkQuWNCfPoG7As1glGV2p
L77C2Nwl3KcWG3RSM8WRIkgcmkcLMPy5H8Hg3JobofIR6l6ExRAnu7Jt/6/p5a96T8avba92DSDw
Mfa7cBA1JQreujRLtKkyt10/jfOcSrmL1SSfRVniP7+QufHihIqBCPhF73JVWkiKP/g8O1Hd5KnR
yrx/13LmwnrhG+Y9Y938ZeLX4xCuZnFRguPi5xWQpW3O6Km7ux7ES9raqHvODE73EHWTX2W8dySH
SJ6JSSSiygUBoEtxP9lsjI6bXG3Gl1udP1ySEmOKUOsiAt0QGUb/VBGV/QdG9LYchXn3+q8HMWPH
DNu23Y3mlAipDX95uaRjwb6o5XRs1uvz0t1f33jECWxZ6+2DMYc6ERUspLJ9/hdku0oX98UEO4HB
jb0r8wQI82+ELhftaKTzPaaPpMWPBnJsfZweCODsBOMRW+I/p2jKbSRT1awB5+I0l5BVCbqQUv8j
B7DrQtpr3o5Tr+dL20cg0Loq7Vn07T4PRNV+mmQlM/yP9yW11vLoplL4CUvXB3wc4+NfPcge0oN+
8xModR+LmYbYuguQG9ZUGCnpVKQZzfNhKJI4rdlsmVHEdML8lEUnwf512NFnU+PjTmivky5Xv000
ykXFAF4oZJJyI/QJyVmofeBFCo2M+iai0n3MII7dByfLVHUwVpdSVfhKYxdKGV0r59p70fAOYwfl
0KaKrM4PLMzmJ3ipiz9dTpnd04haTQQ39qLhldzETFQQ/RuzVuAP8r9MWaMA//s/0khg/nY8kKHr
9N3myKmwank/Mkbz+Kz4HVlSzleQwMbWwvbz45GUHD4JsKpxujTDSI3YhZOd8DM0+cLfTdVlr9NZ
2C9sePp4jNV9Lj7t21KFd2sjpszt03bYA1gkmte9b+DqIL9CHCt+67UfTIURq9zUBPkveXWs8o1q
MWt6FXy+2mW6SUeyQucm9jDwkAft4/vQ9g+RRD7OmvqJ121dK7i1pKXsMATF8GmPI9Vpzobl7GDB
6YdM8kqtyC0dYO9TwbAoW+HFIX5r6kATC9F8AbfWFIn8r99RUjWquMu2fE8SGpMb6wSCS8KkHm/L
NRHi8IcWbbwl5wBKiD5D41I7Eu2LSyMrLeArovTPMk432X7q/8BSsZyVuvu3Zk4GS99gNKa0G7tZ
gCKC4S9xV56A+ndXQRC3sntzZRkx51TLhml+cqMIKp/sgqRhXOHSq2Aq3LDOzXhTtIb74QJ2CEHA
CRJhINQVI39bZtnFW64VJpcq0DsOzvMyVu9CbIUiqPqZK1XdpX4wmvqm6k9rLeZQ5OoyIqQKofVq
kiRQB7pQJQS6mFqQRcSJscX/H/AttFD9I8s53sOOVayOOteBScgUK28jLDwuR43yKRYzETu2aqop
0oAsCIYTZFAYBdMKlAIHxaQ+nDvK312IuhJPRIJLFc9SSulZi2LhzYr6Fu0B0rYO8x/k4GNoaSBZ
poHSRtv5BkBJLcdNUfkn8ChUQ2GdWP2jDQRhnI7yc6QmbbGF3wUKtGjVB/ZHP/Tt7/J2bcbuFEHC
DRX93jt9jtadHmdNsvx+f2oqrwwR3h+mhakyVynB5eJ6lGzYE3llKSLo3RksvDHeVqgYDNO55L8Z
CTbVtEFclJNP3o2hze/esUB3KdnSRz5UIm1zq2WX3+V3YfEgbonHQm8Wx3xqWVmXi9hx3uYD73WC
1NO7DXdS1aSsbnhsXxYmYLBztkT9HDp34/Dk4kUyd0Wz6qj4+Qr/HUTu+lWrGYF/dDPk5lyCmwcX
wgoIcygz0PySKHadPf2FPhaF61UpNfah1dvNmEd1JL4TmjwWSpvESQhcGytn60xOV2aDXoheaTL7
Mci6o8M0cC3iDw/Jw2DDNSIGYYCrDLzl+csIYxuQq0/gPuQdDSgbxbud+18vMMxj6m55q/LIwB1V
SRDK5jjjCHXj6NusyxoxNRJMLrxaYLHlGYDRt71Fz2Rfr3WS0WT6BzGsX0k8mmEvbxzWWjslHCbo
TXDOtjmEvZze+LNw5XPM3afR/dkoOd7A+dvUWif9PXEgHxwolvmREfPiFyS1j45Dn8lQ26uNevgx
H2KK3oDjt4Uk4zwbU21xFmgq/e/ltIJC92MilnrQHJgJtkJjH0RgL0D+XKTKyc55qTLxOUtLqY1B
YaRfB8/3ZHn7ZR9qCf4EzmhxrtWWCElk3j+jQEKmdIXinNwskS6VTuHqURs3GXQRIuK0OEt0+ow+
eJ3MmFReKIW/iLTy3H64wqKyl09SZ5zMgajkAqJpgGmUB4Ux9JpTmmbk5Fcth5Fbu5eGJXC+0Q5t
YhzHrVQpQHxOEnlXsZWWM9GGYIMiTGvHGR4+dLV0nHvuyCy7GKRjxUQkVRG7yQ15ylK8qlYSjY4T
KL5S9SqGwFmR1UcrWAS8lSUdS8ZHoT7jU8BfbZcWQP/N0z4fIlZUfhv5Yn6fn3ImX0P4p9ATAuJb
3s8951t5H7Yp7QC/geAy8FrXXvHMUIzQfTwOLdAzkY3ruQ9gaw35/fefVtH0LKbZiOWh/3m8BzlI
+C9VUy80D5iZGzf6o2XKUv/C+Fw3zkh/ipwu78NQvcWhHA/FViCwCBsbzv03syaIWoN5+tPJJkoQ
Zg++tCAuEtOC+7HPDfWmTWlomTuOM5SpWRcQY01Gv23Gyks0lTy+mc9N2et6ToOV7EJSdKuCe3nT
rwVnMxETdrk5tE08sBgzZfikyrIy1BM5TDKXIoz3B10FZM298QeEMJHzvAvLY2iRpRg56JFGwFJ3
PdVEnbmAX0xMTVy+fyD3B7LSaH96WbO8fVoSOkw7RZj1wY8f+Kg6IISNoimiyf/Z7/amp5ES+i+z
0WA90MOPCOt2a1B51BsANzX7VTkMwKeR55dAk5j1jdJsdkPmaYk1lui/YHGDOdxgRuJ2eTZLCOQo
NlskjZp/9ycshL52tMpDMPoVZdnD/Z3s4+J3ym/l4W5y9kkumfrALOuiIHglAaJQT9SwRjdSj61Z
Y5asPdyM7ituefCzBnaGemK+0fm5P+ZvC7LtzJx+Sni7Zg5Aq+G3P2vMnO1MOPSvSUu+WjF36gSJ
1Z/aXc7bUZGW8zHh1DKMYYtx0YkUPRBMQZv1lcUHrX95JJCiL1+if4x82psF19Y9TJOOBUTBkklg
qTDXOqYAYqFAAqeDHU/jZ2rxnk0MQ/iPggNzFb01uqjIUDInJfP3DC49K9/9SHf4AhtsO5xoq83W
iMCpRKU9vuG+23YBE8Q1xjePq9XhUORTyuI00Z5okxJbCPEUl8cmLqrQUFnSnErCLu9LZ6qkkpMc
FkvxzHH1ujq8gUNzpqSK2PYO1uexTgZDiPaSb1BTcxTy8x7mJX0DA/+ZqQN+1TIhALvr+ZblnsQj
zuB4N2oE+oPo2SFfo+tjiGvmTezyyvU6WtJcvpfqlnPR0/+OR3czNnoYVfWUrUuzdvvq6upFVI4Y
hp3w7qnGtT4VIPZftexySwkA44SaAkqDcon7GNXhboYa4urAT8N1KgNKRQR/UJ9b3C2w6HBkTmf/
nkgfRv5enJIANMcV1uq2evohHU5SdYfdyr5vXsuAlUrol5iEfUD2Q0088zIEnVtHf/qvxrUFXJLg
5lLkK+Ap3vhqd08ZW9X59aWV0I5P46Tl9jun5uklR88OSXy+ktfVuj2TLfCkTIsMol5wOWAomKHw
yHF2/qCS78+qDQN9zhK0kvsA/igcEkxjAnfawyC8PXM04jeeHMxN8WFwDfMpMt8XYdlhWITgQS9K
9NI/44QSBQNiGv3ofXA6VoibHXM90QKDQacwnxo17ELMv0lh9iE+3l0Vw0uuHTdIDbLjNhjBdYs7
CNzFOK5wJZ2ZK/OnVkhpOo3zdPybYOmw1AkTZCTC1Lw9ZzE0LnjUD0UMrmrlhVqxPRqP0EB3dYPz
uW8rkDosFUuk1JqFaoMuPX5/vPFMZbObN3HSXxFDLOUhZNIjO4Rs3CoxrDgQQOYwr6xEaLj04XgQ
XIWGHqWrirG8SCve/eBwO0qDMPC4mwAKbgG8RptK8t3UYsukGjOQ9ZidoKMBH9quwzChs+zeThl0
8SsDuCynguwzLRpjUq/hLoD8iZBKpmjeRleFlEBQcBbat71dMph2vK95Ea1Y7BGjxG0maVS0uNkU
9LJhc8r4I9Bm8rvIKWQ53DAuCE0dqZlhLF53y6km8Ig96+x6Y96u1fwYNWouDEiQZD2b3o6k2ol3
ZsvwlNCEWz6tYLwX0kDW07xd0mFvPIxdtYQ/b/MNNB0EWcO4lGRsuHZsmuta3rKwn6dor9FiRN6m
4jT75fjbRamP+MMYKaCRgieoBhg8IVt0fDCg+1D4d1LQy5s8TSEGj55cyTTAgqIT0OmQTLCdm3Cv
JPF+NC9WbQZwpzJNv8WAqW/lrTOWVN16I+nuK7eGH4qg2RjIXQfvqfc7vrDelwiL3Vni7LoYXUvl
FcQxuMN47knGkPH+7BcfMAw8XWkgSiZeUO7vfQY4yK3KqOa26ZtfIIoH3ZxCSv5aoCnlFhb+30mo
kekfsf2DP5raUvFLCsskJGQVvsLsvo/4wxL4+q8Pkh1PnMG+pAJA4+vczZjnRAUhTMjw0Ek8Zd23
qK7F5m2PFTqwqnPw7TejU+9Xh2+njPE1dKeLGtwT3eHclMkdYB9M1m10i/ZcEz9M1x1gF2B/AH5c
iBD89rOm0VLhIZCkSprxKVu5NVeJc+Igi9htlsfeaXSgn14zfAn4XMrOoox/JbAMrPmprZ5aQmI8
Y5Gl0LwM0FtdtWXRCSOBxptUAAIqdObMZOmZ6IoMsj71qdqdPUET3v7IoUW3/t51vaagR+Q3P4A9
eNkkK1sxmJMr/tWTr+LsHfqqxgZKJTgfRHtUNHUx7nn1KojpZ7fuZK+p14ZLi1vIB+W8aLQLpXMr
+2m4JUubksUYVxaVLopcJiusUO84imW8heiyvs2Y3h9N00zwjPtC5XWVpY/m25zWYPuKJLtwjW6H
tJ0mXqK5RMCcLKjaGR2N54+nshqjpZLut9glci21hCKCt+o1ulb46a3bHC9Wdk7o4d67QKyuTgLs
gNR2z8tbt6kpCW35asBwCYOliqe2jrT2cWgm6fSM6/5xkveYIw0soNX5Trvb6cyKKSXy8s8nuLNJ
LCI/Bq/rfhJFiAdvWKfSYHhdz5MQkV/j4lvYiQXdcFsHjnnEyU0yVuzWO1XuackePl7qgIfk4wex
DqkNqxXo8GbzPHqg+VpjI0Yaqieg9uPJ4/o1hfIXTymbU1E/t/wXfM9KvXYL8Wls93i7fxNi5s/k
ioSxQDeV4SlXE3v/z6I1L2TaYCRffP+A8R721G1SkW0Zln4KmIhsmliZwaaHJw+i24EI89D4v1IZ
eO6ZFHESfv0aONdAtEiGISmNXljTYaSEWW7qAP2KfRqcTUaPpyKsB8TK+FuqY/l45iniXnLJRhb4
/I7crn3jilSmpJN9cRe3FGaJxO2fAbFKRvtZ2q0npV5LX/vAuStme5X4CKiYRQz7ROBaTc8XJizy
dk0bTJ756ufnt9z3bCkOVJlnoZBKOYOU+Oyejp4WCDpTjuW5olAMpGvlKZT5nFlujRVEsWwa+RhK
QvaS76snScLKDx98vWljy3Lc38dkrbgZ0Nya6vREG8FRh71ZfFX8Qt3A9RDxtdr2l6ftfuBwZemb
HwNHyO0KnEq9lZ9eG8Emu7z5zHUQ+bv30s8vS6ZtTf6uOxC4q7YIKZ0z8ncg2RFj7Pk9stRB2vT4
jOx5OvDUH3dOHKCGA095aaJPLnb5TBGJwCjMXQlmznPnC199VNIm3OEO9kibnQuFEsYdzlo9egez
vk1oaFZlpToTOVF1QSnae93A+SN3pXJF5ghMHRzHyOJKeklOx0/1Vwj5pPLab4kDNzTYBOWYUGkr
krv1+BkWMLrbM2EcI1Zr1cqCKpMK9F8/spJWDyYeD6a0pqyY0+WrYL04xQGxLaDJ13RkqsjrcR4y
MuhipE04UaI5IgWv+yaXEDE+OWKdHJHBp7qdxHmSv0OXRNTWD27OJhbwTMgbyMh7kVimyL3kg1xI
0AJ/lY0n4qHZMJh9qWRponzIx1mcjLyqRcv1YruHT1r7QKQgP9UWo9u2XIE9F+bwrKw2196AGe3H
K9r059mbFu6+412bkJuywnIskAYpgpEWZGHnhSDaecy80onuWIHFN/W+q1a2BPVZRPCwi/oR4VNY
vXtwEn82e/OK+09PIyyWtZm5tmnleFq+14AaAjVUDZoaiTgQjvewb+ESjd3UD23Pxy7Ec8vHAYld
81X/BKKIRrQQNrXkrs4wQ9UyUt03YomB2EuY0IWIqkAcHkHueG2AOqLTJYuGlZIE6cBlMtGP0sDa
++/92PJ6d+Xrb5JSft+8F3D1bZ3YbJiAwRvGAGS6H1wRv46Z+2hA9qTyKWbkGRCE/56ANavubBYh
bCHlPRiiSV+nhwUKkG9ZlOlAwtkmUoI9p5TV2N8k8GU+xkVKu3PCPX7QydqfExHgh75dh0ldZ/Le
MH8TeF7p7784QSM6Ec140BZS2QWCpPyRDb1jJmukTjXssoP1nPQtAv6Js/3D5JIQATIvKZ0W82tm
7ii3rxFVNhO4rDx+CvNrjSCcgJApWy5yZkdyto9TpnoB4SR1NTHIZfAdAOeMiT/7/f/Id8zYpf/0
p4TqYsAoYsQDFhpLVPkQKjcHQ+MAyLmm/Z3J9clJO8X0v7sfScw7sxHxS8POUuM5at9D/E2obDYv
AX+BP9uUg20zXsaHLdhzJdIE5VLSadeBq3v7NNAzdaHBE03B3WgS20V5n6h4EFtnu1nS1i2ExsRz
o+zvIL3vJuLjDhgFgGm3X3A8OAilA4mf1MLElDajlnxPCU73yfKBvqkhLjM9W8dtjGJj0fB4Jtdz
FE9NnKUjEt3XPef9uA/9wA40ibSBD7b//4xwfH6rsw0BEdn2Ed+V0Ol/05OEm9qvJzVVLgFJ11XE
Ne4L6iLHaOw5VcWqU8yQoN+QOzvGc4NqPTd12vO6m9l+RlMLgXnefDEzv6br5juGDOD+ORgLWCON
hJNNJzSGJLwU9Cbb6L74BQ1SvcPb7LJS1Dix2XFvsGlbWE4nhwx9vCYhJPniXkZtb1s2NS2wwMU7
/ckhEadkbE37D+qnS3Kmj2aAzhb2ceyLVqkjfhCy05YoVbXLKzL6rwRx6gZV9yqZtkF68DnmU8IP
f6qArvH7dRMSZyUGroewPwQQTyJMn1sXqYASKe8r8bzEmL8ZOt0uPggXLFfd+adCA5Khl7IbecZO
ka3mkYgVLbwPkhZK1xasxziGaCaOdVgSZdWPuYiQAThGyn31U7a/IqKLYg28q76xXvqRHs0JbfJw
W5Zj0zBK3npwwv/dQxpMT5UHfZ0eoSOk7WFWFVvwgenV0TvuE7a42HopGR7S1HH1BXMYVrGE5q5L
9iDvxrwFFYqtqOV/4svwaOavcOo196np0WtF8QNEBKdkuj7FzDJgxmmSGJ9RquXL6at+82wJbNvX
/fqUYPb/Bl2NC8arnkQ4DZ6SpNIFloUH7Qk3R2QzLqiNABZ69BXM+QwanCToISe1TDgAJ6RJrqaX
OXcqdzs2fwAhXdqG3jdptyAQwmR4iurumJuU+TvK2J24uFaQ0nZdxIya85U5gO+OFjaBk2ieYvht
xi2bsxOW6WWqyck2D42qzVqrHiEu2VEkY65/DVeAvFFhmmTGg98CKHmuZLk6x/Tto1B4uhPfIUil
DrF2RBJ2DIiUcmuKUKMvwon7634PHEtIbbegXRLhHsNE+NhAqQibiOqtDc6GS5ixKaLFhBytGI7u
f1QBj3JELJWTV5GvLhO5sjmdcZGxqp4yZ2YBX8yPQQYZmLN9YpRRKOVB45tYe/XSWbiE1ArtY7qH
d20wB6yDCkgDQwU7MNDponbkyE2MTNrfX5Rw11dAGptMKiWBIOJzoBrMTcOApORRcvRLKE5N5O1S
hMQ2Rfp0cSDcRx+GwLxNZSLcliAk41y1dxZPtd1y13V44/7bwbQETJa+OfyEIwmIe7qULKkWpK6L
DUnF4/0GJvDyZdcH5MZCkN4xq7x3YtXtEmFgBt8JCE3JXME1k13iCP4+EFf/HPf1fvBTTMDAj4+J
7hGT+K+9dQr2DL7vdL3rIypYuTCE4fMXp3L1i9LUdeJsornuocV0uwtcn3xcI/1GYaCQPh0NbxyN
hbS6dhwJJve20QMs4n2FYHPl53REJlPTXzBEjMreH7ZlPrGVGKZXIES1p0ZBGgcKz5LLoGj0D/hX
irQEJ2/i54Kpa0k/C7l2M4yccM48vRFGjefzUOHAKOM79OWAJJyV1uUaUiolKB0+jWGqtlpLC4mF
xrxeWPUXQaZAen3Ldz0FsI3n9DPLbLCb644MU+xbT84FqyYv04bkhmAd5jj0HtrrCKFkOYcSTcoU
67FxZNEKryvZYhzA1F/RKV/qqAUPcO3KNd7PJcgFPZsbY83cvwULaEpjscsnHYTuig+H7ZuYys2f
7bdz7g2OQOtM2IrLlrkzbbMQ4kSt9Jf9yszt7o/rVtmkp34EcDkirp+lWruercLBnmzFZrzF5TR4
CNp5ORh9ChqoiXX3nCoKiGo6OvpW8MAH55L4t7NbBYSiME0wuTKSDVqUgVd7Ylp+dUr3bwwMjrCJ
K2ghg1yf9RbihRV35XE1qZjr6fppU7yA/7Iy/dkT6m4jezFGLgjke4HL3+hYFJ5zJLsnWos/Pa+4
LzSFPtyR8By99coXARf3kQmRqvKejmrnvXDJueoHVE8NbgHXpqAlHiwkfFi0nBt6VIErp+2U/rBR
yTy9Xe5jjRqUxfQJJwqzZaG+zyOlnHk3CAQGGL3P9JhIKZ5IQ+gPXDjjNeUSTkXpccGJjnpOTQ02
ore1OwXRQLzDVuC0TKxNWillcqtPbaCJTiGFTb1TUDGmGAjL3qzg/ZWomTC20/VZX9MMpbpsVf9X
KxwKkj+LQc6ikCsrzlnPQcRoRD/qHcsu8UOargFHw8QRHuK4V7LqckghJki7fW/0gACB63r96+bs
Nb5ffrYblO0S7YoFZGUyBqRAsekgUkedbW5yc8+z0zfi8VCBfZD8nVJlQRQfDXbsUubWtBkUYBWZ
bw/QQr7i2wQzb6AXftxHm/rDyYOQQH+lcFFN9ISpE9aEYyp9wdrD5HQx5MK9smVrauLtPDNAV00Z
DEN1meKstY7musdR+c+SLdbwqhGfizMFFO1CPm5dqMPf+w8Jmileq9un1E32CPT9tFmTCIRT0BzT
0mEPwyZbA+PMrIn7Wlm/QVgs+hrFZJ78Uy+fYWhnW5XC6Z2x4dumMwbExMi4nF7PaHnFoRVfC/wl
nOMbCl4g8XIo5Tau8GHtZUjISW2eZeJkLA3S4598rTSGfqRkoo8MmxX9kbGxuJTTn9vVdPyDojz8
cyn8OlVbqNgxXQF8MD1sW+LidWw1UjbqCM7TQECjWkpPSQmSxqi4AcY08VOHGYUM4YQBsNOsotLH
8V8D/aIlZVL5teZoXW1wHiH/13WjkiJABFut4eJdkBdowRRWr6L5z8iczNsytnzxWQm1+VP2TCQt
/kqEe13Ds14+zMDpwsB/dmcyf1E+XEV3Zr6SW2NkJF6PX//1KEossWuQsnqHlmgw5Oi5105bce6c
eAnLTBSGg8n7oJeLZANg7+DJBuQJisTt/DigvCAbdXy2q5LfY9Ys7EAcYuuNT/mg0opIG8cvOIlU
09TmqaJ0HdFa9ydGjtcQ+lSqJd1/CugxxdEw5UIqVOECsGT7JuFvp53/guyWq89XWbo1IOHy1eXH
5St5aJBG1OlZ3kPmkhklqhBlclV9TOAzUko0fYvQyRW49uE64bh3TZhNycZlQFpo7QEXp8QmTCkP
rv5BsPqzjCVlCRbdOLBgFACqOgt5rRSLyTbpjmw4S6ApwXHMdEylmzDx1lFOQL6KBSFp562AyGRd
gRWFAT2gX/wkMtf4Xx8XJfAMIMXjCciBHi2I6balHx6Kqzj/jyxuWDbyiWnZR7AUsvVKQ74Txi3T
benl16BzRYXAJpLEMvquCFlfB8FnkjEJ8rZilZqzB8XTqOxqCntVQVFnTeoWI+D2u/tF/6mkJ2xt
s6YPEXPakgZnw0qb5WxO+ZpfaFUWGkXd5OmC1pWLH5OyMojnTLN0v0RwpRGIrzj59inZzHzYaHTl
6xJNc2n4aT1MlAcP0CpEudUu59HrvtS7tMs2mvIink1Rclr2PyE75+OayXJlF7hz1+Y83k2gj5xA
UddXWkhIYroqUEyRO43VgPwqCFrYUG1BYyW0DcYDN5NORIAg7J/YivEdzT5jjQuuGERAeWb4PsMo
SW7qrMkkUp5biNcHoQe0bjw9fJDHXKQtkmeQXF24C+2zO32NkOudPZ4y2/3yBlvGgU/ffBJmP8QJ
c0+3WFeQRnqbYvbTGoqvzjedIfYzHkiJGWmAgusBrd3smQWZjqJ8Q1I55EzZmo5A9mSznl4t1auG
+/GE66o8QRuxukonUVH2XDWNBWZGcuCjJC7a/p2BPG9k4iwL6vEPYPRoA///0e9Q3Kaj4OzGiACn
ecI9Mo1Qnci8i7xEorBhYUld54+EvM/ALuALQiaBmFjEm/iuXM0WLlQkqMI1tfqR+jaV1UxwT/xA
b36t7a2445A/JClAkiF1hv5KAkO+0EinXNLyIc8/26KYQGSPbzUM5r96NqCsoYk5Q/8dcV1Svfm/
ET0zc72gM61n2CQwbdnDPYt6xg6Xz4x7QVDju4t3jvgKDTwiLkkfjemcG4ZPipFt8T4R4JtRBaib
kvH8h/2uY0te7X/1dNV/jywqwQspjFcBSpev1KEqc/4VZRhgfi/sSumj7LQNoqiV2qH5wMok140+
TnKhEfeqNulaTcJ0fKN+JgDCan2FRYo2vA4d3UD+6zXjfpkQZCBwzane2qjwyHTu9ipwYEHkKnTL
ElwVlK26VraXZGz2s3/sfwa+6VOooLBgCTzLYgVMlDAG4hkx5k/cRemabq4fNrToIiYE+ZdqxpfX
CSjvXbXhXnqnfZN3wJaUW6A9FiEyrSv6cLdLr2rNn1sPfJ97w/oCIoip2eqDXmD1tXFXcri/MBn7
Au/n0Dh+PGiDYNnBozSRBVC2cJtRb+T28PSFHWjDVxr45H9ROlS5/ktS3OivmdEB7n4H8hbpux1b
5P8pPhTc+3U8rW9W7WMWATEJDnRChBMObQNk7CMUQ79cLb2Jx/X2SFuMJaZuoSacwm6gGT0xZJSt
a5RUJhy+NR9j0RxYbBl/2sfLT02ZvTipnsGY79s5uA3DthjcXouFmP9DtwWAfOyWejtzwW1NBMFa
RrAZYKmAKRtSf5e45l0CJ8G5vQV3Fjx2yrrWhnoPjbDEmoGaRT8mNMnZ8knQZ6lJ2+HY2ASqjsTg
U2qQrSTFuI7E/DlqQwbLMrZY08S7c+IWajkPScV5wFEjIEeIfIeInU1MQfGYdcBAIqQH2NEeGiei
l9zN3JNvTZvsEdiYiER+RNq7ccuW3KMf92SwrGcq+0PPzMmudyw4dwDxzTsGkxQKUSKnJacCFJI3
A7ivXLXSetkkug1mHepaPr/TtSSJpu6Xg++hfQpxRarKM0Ua2xnBfeu0o2/r2xFjG1vOZ2Rcosh8
QI8OxjgCa9xX6B3ThbhX+LN5MDKlxRKcdpFcW6o8QVu3W9Qo7pspqsRimZhZ7JEzGsIEePfdCQk8
TDF07crsopGf78E5YRuvWXP9I5Iw22U+ySJXwvqvRgkC86VyLqNXMGum+G9/Q8GnA2hZDd9Gy8SP
kUe/qI2Ob7DRNf1Q0L7YbatmllFabpTkHdpeWYAyk/AwdfRDFVY24SMEKAGx4WVCecTyjxhcFvNe
JTSj+uOBXt8PP2pZtU6Y8fH1pDI6puHFOmklxuKqZifNGQW1sg9laFlvhXaClljmrGXrKBT4Qq2X
vVWLXUq+5yOFDFGARPI0GNN4J26PRejVZZcFy5XixfhUPLyoCC2PEEcu3P4JDwDOeeNw2mOCFLY7
g3b10g6RHh4hJl1fKqgg921PL/TMgEWPGzcxuzgMD7p2mlziSmPOHEus+g7mQqCz65ufDS2P4DN7
HO+FKNUTLVvwRoVNyDsLib/RJbdJK6D92NMso0GhWHSfFiwXIQKES7sgW8mnHSm3QJTaQuFok2uQ
EzLneQTS1n7abOAltorWWqioBDvmXbGiVu/fydk7lYL+T8jlLg3FOzwzuwZxHtbDqAZmNnvGrqAH
MurjtZ3sfiucv8DuN8JqkZyeUsRn8ZoJIGoD/VMjDgMbnXv4F3F5C0yhM4favfjZ+etpTehX4nVO
8MP8N7o9A/ARCM2kOeXvZBmMK2ugnwnbOMp9zDh/SRoYJxHut5Z2SgmRIcBKnVgXSkDGPrNehXGd
QKNg5bf3PBL1AlZdXynQOxM0pcsiDTk0QoDLy1a40Ix4pC1/LLqcSIxCTSd7qQkg2cgxNUV+vpJc
8QFrVDfRRls6UBt8pYSOIENRegUOFtBbYY+B7pgQtj1RxQVjXwckqgAR7RddMQ1Z9lCxYplvuI/i
vf0d8Vc94bbVMuAn7HNbdpZnV8zcJFbssPZxu+GQdpmA10oOnfFLO2iQQbkAOGv0HFsmg/KaJ+mE
2CnicynbCzhrjIS4rqiFMjbHGlfLTqCMUXxMwBIHz7b6rgPH8OiTWcIQvFcnYrLpMBn6swNoHD4j
7LR2eG8ffj9zCIH5mDocL0Ob/KNBcNgXy7l4+/aYNyaCfXfq+0qYlTCfgFbx0NsMUuLdvh7WsmG2
OG0pag6Qzv5vAvV8o0hz0XAr0F/0h2CBU8qELENvZmDWW5LmxhH5Zt31DvoTwg6ZC4h6wpWZys17
r6ND7ytYEqH0X4CMg/B7wKdy8x9YtnVf3oOyD/31YRjjkwwMuvQ21A+7t3tHCdZ0ip0XYkSv1LWA
SHTK4mm9H0rsGDYhdeqioR6afXz54wHqECEpS3HVtn1DWqC/rPR/XPgaKLRBi3S7ZIz5neVpZUkw
SSlekte5REb4hBHY3+q//9sHbD8rWCZvBc5I0/UcyGUwUHiMYAF/qq0v4J32dwytW8eld3ljZLdR
sNLN8JswqIOwApZ53zMT9pEov2eR20M2fUssPkqtDj9Hb1XRhsjpXnkKD95KhtGrAD++ur5eXuk3
R7PQBehzyNh5b/7H5lwCLaKq5TFSlgFPKk0Ka6DWqmqGLGj0/LwT5dBa+cSqTfGm3agwfELNV5bx
xKO4U/lXOWYFMId/qwzD1TT7G1XD9pf2rKgaZieCJ3Ommj59iHaGnbtOXsdbeVcXiDYQIyVQnfiV
Ku5vwcSw66agTEH/nfxIqhWlTShGWjjsisKy9FHXHLIO4+fAyOhKZOF3b2b99iNjo9Ejrk/rgCy3
aGeD9GTUUxy3JZdywCL0CcRmEq75zuAh7ARS2AKkZM8MPlwvkVpg1Iu2PTVhDgak8mdm1PvktW6O
jCxvCOO8N+JBV/3gRzNHwwF0gxWV8f9FZZBmNRZZMiryhqvdkq9Ck0oCZugl4sR/Knv8fYz9JSSm
Gkd/aa2N/ggwkKsuBYfTb3SN0G9ff43WdiJFprFNvQ7iSx6S6R+wc0x68leJ8JDkdgZ+Gh9l4cKL
D+LaKy1tn16/QN96I04RdOSBPvaF9/5n72kMRu1GTpJq62YX8WsYQ1kWgefMArdL/g0uUEdbNKfL
+4opgNE9EHPaOPpoiQGfOwjxFVpe2qGCd1pOYyl8f0kwHFVc4kcmCh8ON7053TuOPFXuYck9NBAi
k7hTjDy4mQduYcbA+bQNLnFTwr2bX2KroVQ2MzWzIIXoKNaPV2oJzuM8Z+irz4ts5qUN3EgaDlWC
TiCGP5hK2uedcolm0ksZR5K2DqRtrD0mp1K8zFm5UNmRShMIxHt2ca0niVuxy/pIeMTu3uHLdkr6
OXym/CYyTY/3MCP4VptdN4eW5AVpOuD7Ao/H16QPpj3cPOnVYf6lcC3RVQD24LVGZ8w7VldhQ4ww
cezsLe9oD/QdIRRHP7racDai3SMnyZzaQvV/AL/tLN9Ottw+bCnHrxdRRXkgRicudjCknXDTikEx
az5FTo0WkW9JXY4i+GsUN7qs4MqfHkx/LACacgyZ4tJJyvVYKMKzq0MO8b/P8qXeIVym9zIRmaAI
VO2q/paOzMa56fvCAJCGZSbj8GYBFCqKNvW7cY3GXloUXWJJzmZORHzKiB3DD9S3JF4CVxwMOBJ4
fxCTJWX4rGear9Mmy0hVzrove2N2PP4ToiYnzCpJpGQMB+YZEfxC5j8eVGQ9D/5Kq7jduXAdDHOw
B7/GYQPMn4YKl1ot5CTwWohlIhgwWdw2SBKxDLS4jhHPODqglRSveU18c6+7yMEnYWgz9bCqDXYx
eoX3BV5b95Qdv7j38JO2+soGi6K7ospwADIxuDU2aX3hH4HzohJF4KwRsq8FXm5N5s9hRlzEIXVd
aDkr3oFTQKo/LnLX5Cni0XIaCJ51EkleGQgRJlmT+UG2WU9pixt9nb8PIiSQ+RHc9Y3oo8eJc+12
HheNqpVhZSx6pMFI1W9g0m4Ozz793djmWqUsrbTHMpKFkTULWOUW2bck98kizZM548+we2ph/x+s
mqnZNPtc2SM8bab0qPlCceQAooTdbO1ASLYEQEMZs4L4x+V0UiVTfa6w59qFS0wiqVPxS3m6DOly
YI3V8/Qje8x5eMcpsuv3F7jsjLr0u15sLAw/K16lZF+sJvFqMZZICn9MTLSiZwM/T0hCx7La5xYd
rvZoMqQRESCuBo48kDwEpXO868oZBb7Bh4d5jJXsjXd53eg6q8w6Pd4lTeLzaAvB1j1x/JA0S2io
1ahDngvLnKOlGw4g0v/BZbjCcauxwFyxWZobLDXEgZiLT3nVPDtJWgkbhgQxzC3dLOTR1+YiX0aF
K8NMqKvxjMFC57vAoNMlU5H/8bQvyi7DWuGI3mQe3A2bEWlZgWiLz2l/P57FjPkC9JJC2U39tJrE
/LCzMYUNQcz3ohtyGkd6FxtgHgNyK7ejdT6N78X+1SCOukeoO069oLbbCZ+PpwTOdAYdaH3JLKhw
6JlOPZNu3ejJ6AFugicqEVKNpofNcQdLWnWj2M0RddYcMq6rAF5JITy/uyiZSgSRpmX2TtA2I6Ie
cZRrEpeNTdB8bmn1DSSzKyBpfL5sIei6eV5YwsQMY/etmMWAjrgALBKzOYAYDd+9x4a/IYBOxYof
ol1Ykx7Gr/VXoCKa9nhy+YUWXl2S4eHPkBUJODfBS01Fs41m0lyB/jzFlrv6Jj4KdvNi8PGR0xL3
mX0oQfy0L4iq5f2gM/ZiAwclenyqViZw0PbUPYMrqssfoXvo/fWuzbQuhZ3qhTYEIxvRguZkygUd
UUdK0xs/8/PfsZcgcpu5DSx2ZpTQBvxfPhWtx0SyRjQvNE4IiNP4izv6ieuZp/5HSSJTwBFCSjm1
rHS4HD3pbZ11Uj2NOO81vYKLRIH9idOZB9U33RUBL4QXPmwsXWMMTzTbRi74RKsI2F4SemLbe6Yw
QO8ukGEgHi7UYWZroaS1KsB5BVFIr2B4Q2j9BRCgojTh9CYg2HD/1TFE43rUEBtl+uoR06jsWAwX
PPdRvxwrqXJxcq06SG6WVzTtM4yid3lmfY/Jg9olQjjB5Va9rVPSD4lcun131Q5tTkWZ6Fc2kjN+
aTisgWMqIn0UysJyerDcmsbjYA+ebePDsCW8DrdKDD4kIQAvWhSRFxmWnRET3e20gWsBy6gq6JiA
DMWH5jBTQmb+ZlP+h/aCRUsHilCJhkHsYhEfrmY3PwQSWvUNJBnqsMCoqI/R4VfB60zKcsMtsNK1
XoHqv38DOMJvD74xzxBLeXlOJfYyxfZT6+KdJuj9IE97N7VxHMzbPRdWtxNJ6IiqVQmC4PN+Zgh9
trfQBwut8F45ldUUj3pfvt8fnHQ41i00kFiU6PoK/6mj8TN2VBqd588O+AJ6ZD4lbhgyKjkdlJ5+
+aX0Awjt0+PGI4mScCCgAJLKh2ml7YwxgHae1EsxdJntJYeNvkI6shHKn/xNXwzReW0ENrE6OF9s
kmU1Fv96IBJTOQaV2j/MgKGgNs5Kf/x+YB3oF7V1u4SwbIMs6hyR0SExICTMutEkaEtpvy1TtetI
WGew9ZAvOho4EM6WhUP1n5p8VuG0Ph6sE1j72qxD3lxuaPmGB5qsuqIO8dyZSfdrZFQkzyIs+A4r
bmkSUzt45ZsEW3fxGozhwO1+7OtpxJ9da09SWWUZn1tZhJdRX+8ilbOXWTuZvo/uWcysJKYSMVZT
Hg1vsm/iYgaRpDSqLOFfOMhFgEzZUrVQGaiCTxNq9i2y6V9uXwuD4ph2mQvFvXK5ohsPqODdCHCx
StMuyedQpVXi6YFrMCI54PGRdV4vx51ZWcvfo051SCUxJYCV5PZ+7xpm1SDDeMDdbJKLxmBVSo3J
cp7KoJ+uBfsZkUI8I5FDuFq+C1dpHSRiH0LlVBjmWZcEYfUve+nbRwK/eKEHmJpzodRnIJbj7epg
+bXaDsjxaV/B662+9mVyAMyrdcxDdKlhJeP5vsadJVD1kQLh8/UfNjxV0LX9vUt4phWZpmF9JGvB
i7LS4sK8/zDAnMkLaAXxdP/b0OvEa8rEakBkvUCUewJDFjh3+kTzVok3vaMzn/AG1QytxJqSnFOr
myoK0G2TB8CRxKlKaOwBT93iYsl6btYa27vkUb/kIUcn1pTO/jK6gEeBXmAmhjKv8LbY1/9FUJ1y
sk2XJuY/VO3fLT/PqQFQxeJit7irJTVzNpv2pMyKxv8bdpT8W1a9G0LRJlRjb03qrPsqS1spOG6z
G9L2Hb28QhI8VzezIYu6MgebZTE04ulgFbQ8qfc3TeIqmgVACosRg/2bZeLMpez5Enf4Fk6wJm/j
Hk4BLb1RHmVlHEF0DhnkSvuVWGpexNU2OH4740ROpCMPiLcOy+qdxND9Yv9THbWS9qb2iP/SwisE
FKH7cZMPXyGCcGheQaJRWd3Jw2//Cav/SG9AKeC615tlIU16yMrSfX8ExBZ4fCb3il4UQ8uNZ1rZ
NdT/5Bv8Tiy9yE1sOi9QpbGgGfaigjGa0FeiyqPeW/DxYY3O4675OvkjQqVJfU7EJMVTrhzIZsrk
1wG8NP0W2jPCf/8CLCUPEkCGe3wxBXC35nX59asnGfFAlNSToEgLef8+z2o1M90+GltE3VFy7uVe
tWfg44PTvBfwdJog0PDfKMwxlSi22szDTiTsLXkuZqLOwuhYVDUd8jNgFZcFZhvgNlKVkP9E61OF
+Qq7+TvtEUbs25SMC8fL0n/yQrLKqFBOhUGxbB5Zka3Bt/z7Lp6ChG0NuQFo+XErqld8QaYOgioT
+Xa0MYUlnCrJ8dyLpBX5Lef6hymVMZxpdLyxOaC7GU7NCQnCgStnZDPlRv3Log3KBzNrdC/ijZzy
5jVhCFXVX7GREzfZyP9GY6/XlV3JCv5Eb6n15iYIKU1KB2Wt6aHC5SRQekPzq1jDRvZPxFcIrQLG
9Ye55bdPZlJB9sJCek6pPDWjxHSZpKdGlVifhiyuDEhnz4gMQWeFkIPgemVSwQWkVDSYCdCm7UeZ
YE18xiaXhMO0f/L7G2MrmaeGpF/Lomh5bY0sVFWYX7WL+RNKMYom6gscsYTcJcvpmPPmwN9iyiOZ
o8v8nt0J1uSu9kNyuf6kUTnEZu13zDHwtfo+EucwqwnU2CONsnQtdHBoX3pldYH8VxKwFLLaYK79
z4e3y4vsqDc1ah0W4m0PeHsIbsu5ITu7NrqTv2SS2hZYB/o1rrpEC0EsL9si+Km7AS4BJqjTWXq9
h2zn1auYUGEUtmOXZclL+QK4y6cuB0q+mlSlY39QJ26/uLd/42MjdRNoo2clG1i/W6hKxUbzh9n1
mSqDqlbk8mMtmcD+S0/xHiWGvkoMy0mtZnJnBPaiA0CgmTGWIVa8MbN6BZsoruS6cRWpZrPPUytu
hacfMVDt2YG7yxlXU/pfxyN9RL5Bo50AWsI+8nK/8mkhXTk5anLf4e9g+wrsmsNKQUiIqazZ5NQN
QSO1mcd6CrEuIJOJMvxJXN+G+3jWdU6jLMAblT1ujN9xoijxYd8RNz7dJktyXEzr+TU/AdBSWPvh
McFw+VqB/LAfambSK/K6jPIYV25kXMUXEczcwk2ySjJ+7bTUMEFUnyHVSk+Glww3iR2th2w8Q/nU
/HHuEqOHmBqbB3WEK2cphrKquvLvnun74LDKfy7PaO8NrS45h12o9ob6jDbbMwDx9bv2EABsG+JP
aO2hBi6b8el/PYMIsaciQWPTeigf4E6Zri+Qfh6+nV140hLtQKyLs29qmTCD63U3dWgOGaPyeUsR
AQWm+CpjYo0LHx1QxDcpVi6TpbGHtDKkwNWhfoHgKaQYGzA8t7fSKgugDBSMgNGA4KE1Q/9IqDIc
FD1Pc3A3bmTlbtfhmg4TFAkq9BR74MTxJVc5OL8Or0QOq+ukFdzgCPybk965SsFz/i3xkVeM/EcE
K88gwaE+ZeafGMyXYAkLpVkbBytgPYOpPmOtrPGnJDlS0AWACrdKhDE2D1VdrT7h9hi/jhe4EMIj
LqcUZ92fKC9BAlC7C55gk52JwcZFecs8Tg2gf6DA/zAZRAyOJHfZNZ1AfU9luS0qpNkpy7Nch5Oh
QEUbcDHPZDrM6NtQC5LIDxr2pEPyY3cXZc10i973BUclyFBzKpatw779ay+AoB/uZyvP6iyARoc6
TbpovewzLJ6skaoH+l5jTPmcT0qUaG1QHFpOWs4tLhFfoCgqX8WPsLtcyqvAkrWg8f0v1w7Fbyap
TAhodC+onhsYODKD/9NYpZJDvFDVKJVCRvXlajIaQIAf0ibTuiSOekD7rk9pnsyeytEcBsAA+u//
d0oxGT9q7twbsAJiCARXpC82KAZ5QXfn/ntehLVLz2MZ/P9F1EHG152Qlv4T2wRybGyyIMpMn4pD
ZGQyESUUTfrzJTE/EY8PQauEMrbR6m7pRn2Nfs/u8VslvpQG3yasEUyUiZVHnCv3EKRbPRP+R+JY
h5aIlMOdSv2guF3h29IF0vmvH2ATiD87Qr7M16fIv6I73yHxPNSA3C2Jm5ZOlayiHdhRJnN2IG8f
15xJRvy54sLo7WJYv/1pRrHMFaovGZ1/oV8xRwaEJ72IgyyLIZuOr8UZ/7+7/n1K1Z66lDhLfZOC
H0GJKwFGWb/p+4AniKA1JfhV2sj045kA5SqpxdjWctLatvJ8WmaB0JeUBGriIoE8Q0mhctW8iPlw
w1TToYYsvcTjgjXkoKVEBlv1jUgVFUDyiajMLKFovGTzYWAIXI9wKMW03Sb63UISgqq/MxKKfuaD
eqCypGyeA4lHgMWEfjLPqyCB5tZvykwg5IlB/7n2ZE41g4miN9DQ8OiUoLlD9mpf/3R1X6CbJ7N8
Cbr9gBFHbMVSzfUZ1ltCpuSW1Z11lglePjMYu/sd+C97sJCmicxWMMMwj5a3OzzQjALT4Vtr//iS
u1bp1NBYzuGDbf4GKC62WH1E6BuOmpRgLnwKHnVzMT7FVdq5Lw84FRDmPE5/AlUlIfrWmzbUCYjA
mqw9IgDGQAXAfC4mw8rVMNnRHPocByT0xxHeXucKLsH6fy0qpBxCkp+TiJQAacSMvoqhYG4OZq/U
QwaVWl0Qc42mX6TsDtOgU29LyznC8yujlDwg86p04+gLNNY35zgooT7SPLoJDLGwZ1Or5xEPlyYW
HBj/ovAPSI3uHlkIMBSOUnfqxcNc7E9z03rIRtX8pThpaB6XgA69qM38/NU7/54eqdLLbeAsqoFK
CDFKMPxJWoAgOMYtI3q1gwaXnfq9as6eBftcsDaGjYFOVkjF4OWion2EuadoYTe0TIMaX4YtBPwH
WernMWCk/cYezd8E8T6XulSYWCBwshvh9U2x4TiC4lCQjUftAZWREizWi5jFnvTG+zCkiNpHvhph
Y/ZIxtlrM6sQ7typt1oQ7hKxgrjpkc4EjnK3z7YwIqW909X+Uoto8Nd+hCeU54Xh6ESVV5/vx+wF
zT4QiwxMZTFpHAu7Gnc+NCX0qAapTo64/MM+O2/PvhSRSh1123KXrjDAdmZ6oQbJCxrQTCdVdIJi
mUkmDQ5kYghUNl0EZ0K+dTVUhWmtw0XtAPORrjr1VQYESRsQol0ZqyIyTzKQzTMO4QZsziE5SLkX
nOKFUJjYE9ht7a9nsAqNNZoBJXTw5b8/PG4h17v470sB7i7+mgMxz2FIiyybAIsyDyawOc0Wi9bS
WbVhFgq5xBkqEvOdOk5fneavU6K6BJEtl219WYCcAjJmmYVc/4Iy8/d3+iAkY/PRTnFRYAZwKF0B
Jqf2MQJpPoSslH9xoXK0GsjawetjBBPvmBEnz9ZNqAhxHNhyOOH+zuQqKRjCsIEspEKRYfz+7OiH
jeZNTb3WTdW5rw6/I7ydMZLEPGbvNL3SEl+1Cg6RIHL4EzH7N7Bse2DDXgU0JEUkpSHYVmrQ0E3O
rSr8PhkdRPBAAl5RFqBtlQuE+NdjCm9qplQl8PdMqo56zNtH3LOf8myf51gaMeoN2aC4gjzAYTX3
Sxejzf9XYvzeGLk+Siz53TpjtQk+GfqbdHCxvpyEUuCiZql7jEu2uPyY8dJHOwQXjRRnk1+bf5Y2
t29JqwgtlsAow+95Yd4qOPxWZvGoi+2aPS0MyQk51lwoEqPbdF3BgJWOl/Kf/zVX54Zi363Sy76E
EFPwGteHQdJ3YArGbaZMlPUXzMyAU6wY/PaW0lWOdParYFUD0ABz8ercLe6bPvVVIw0VDu5uBM4k
rhWuM7GgBXh5H1ffVgBKEkY7Lv7cGi0mPGrZ7VwxG0JmIElG+VNHkimUq0j3V/FzSiWsEYBTnpJS
LZsTsLFbTqNGRVdxEfqEndFtSke6ZfbIUGWp4biXXgMAU0pP2+pS+ilZIYFf8T3+EKMmDUoAkutJ
GejaOEmCjjJ5XnLqjPdKa7HTzSy4ZfxZiiklWPeHw3KwEWs9gqFi19pZENV/FBdgKXSkFGfUnJ6c
c83H5aTApkfZp3k+3l4WWpyY0L3Qiim+qvXPUwtQdpbViZfPs/SHqFsRADuCMOr0wcCOpdOMdC5T
EgAcnQDgunvAw3TT1w/0OFS1Nq+T/g9g1E69zCLHnlAPZUEg3p6/vJpv1GQ30l2qmXmfsZDFE7MO
myiZYxEZ7EJ5TkSVZNKS78Gl+/0PPQUGX7ont8EHa+MquFebWrK2EEa8YJZl6QohQRmS7FOjI0KB
FSrFnlzOu2PuLJqhpxUKVtcPmZhtUTzWaxA11xC3YaxNTy/bDI1mqJrE+1DrCdeoy2wAvBSjvZkj
8seOTdMkJYkLo3b2nvwiznT1mvn0kTATk9kvMREGc+7t7FPzOl3R3GPm8XGvy7jSmzkba3Yr6FcZ
r3RG1rBQvfEWHg3Im5kZqppyJ7VXlKqJgHFh+VEdlwtNobN5u8TmP/qBAMT+TI5AYUqO4Z/wIauS
IsB22Pekm8jHs1TdOmHr7NVYlCukcLGit5O9mSfxOxmEDuACchDRGBZhmrfGKPSpdN+2OOFf3liy
uVsSaWZk3TrK87i2SfDhs4WkKLt9+RWRT3ESZjWUmTEee5T7TwiJJ8+s44FzOxBNCUD3F9JKsMCc
mYLONW2AiUULlLVDDfmtAFTnGJ4hAusb8SJsHjfbn9DWVtp3qzjD2E1j4wxXIMM6rNlHuR+Hm8IJ
jcvqX/c9Ne+GRbKjZ3lVQpez1+5MEVjFWvqzgQjXKuDrL307HZmUu3M003MbJMyGGKzf61XNxE0L
YmjJvZ3xdb5GGKfLO3hfYd3P0AMDad/aAXh4/ENOW0T9rV81jkuMELtm3KWay+kbtQlIjZL0hyXR
QNHMNNhIwHrMJ2mY+I/88i3ZjTygLk40DvdflknyOYG3KEa1imUHbWmCoIRSoiJ7wlQS1/Y60xXV
uI1UMLGS/EYuZ8/1ZYksnheSMhHWWMCCEZP+ZzH4n0kKFj4AukcRWaIWyKMSTh/9zVIiYuye/02k
Poo41BW6zE00hXn6dYeT93AM2AoT6oZNeOtviwIUSA9yeFHGuSLxq7aYEUD8P9Jc8liyl/hlufuP
QxpuL4wRqtHcDwb47Rpl1u4hxVJJe3+er//zr6USLLSjWK3xoPdkwrySLyszFsYfdfF1pIVMjv8k
aPTyRcWo0urySoEFc9+WKKC5ovUkhTTq9do1wouGYm1fcgErvJyinje1DZ7cCTAvOVPIDs2ErmOr
KoSOUKgwkDnBCcVRte9HeDFiqB2+/2jduTIjkIcB7r6RtzNH8D/R83l6tYx6GNHcrLn9W4bP3SXh
AO1msxpTCUBJ4CY/7kJCPIRFselk1hgJdFN/JptsBFrhffCXDGhFEm1KfWj81tgKojw0hTLBUU8F
kcjh3I47zCpzby3/2EJVh0rZqDlu7cJ0ynU8viksmG2cZ3sEk0MlzroSwnZHQC/cExA1yI+HzSn1
r6lJl+zkTPm/q+hwYSViiWd7NBGAd5V4ECn6OnGox85K1KwzEZJdRxFxORJ6TBG37cCVvRPKwSmv
8VNfxcvg6sXT2AkT8yvdqgilBIXY4cUnNvUlwnCGXQMkSIkGmhi+8XPiKAVr5FC7bCI5b9kXfGXR
bApQvXKG9qMcYPSZiBDedtrk6E2i6U8iX/rAsecq5DeBcDlNKOxPp9Az8wiz+Um4WOPaW9yfkpmn
KYOanV0NYqckfN7+hEEqTC0D6t6Q92nTH/WKwQDsNBliseimXPBXiXcIbj9LKCph8he1b8dsvZVV
1WBGJP0Kcx8m1WksgyItGBzdm4CoZgm+v9v1qYe8rZo2jhO4d/QN0uY1/lYJxxj80UpLjCoxsqfp
fMzEqJ8umWJrX2zJwhOv7wdBeyEAvkC5nLFYsvVkwgBEkjvMveerxTGBMgIu5LwBJ3/5kWKY6nFm
I8teAVWiUkLbDxOg/f94/1Ddfp3m50h6RcSDpbIbd+X6Z2PsE1bHwttHYtuxDWZXNrO39E87yxio
gqmVWBjmBHQ7hq++wYE+CwS9Fp9ANU3gAEyJXDoXDj5axd5czymq4bCrFkFS4y6Po3CHu3WIgdUq
F4hvMPGlU6g+kIykg1YzGF3rTwf9/3S8dErpICiwE1E9IZIf3LGi29XR/pMv5w3rbQ25jfdZ21/K
Bv67fRQ7QNISo0MMTzFeSLNuYrSnTuWPvtR2YR2WnK6w4W1cV20bRJ+/b6yBmq6Fsss42aCgUJTJ
wfGdRoKxCGVLfqR8rgW+9Dnar4nV3DyzH0G68VOs8mODae/cGeMGABG1WiUfbzcM6mRjZxw8/LPM
uychivolmtrHEVTJxD8LQJmB6oovE1OU47LDr/T7eeubvB58Pi5CyPS8EKsSH4X4R14WR9vXy9Kw
es+eYAtP37bNAW1bibgwIsWkSb6AUNltL97wYlR8oiEx0upyGYm2+8EjBZfaTAE1xwImU8ooU/c+
b7CdIj1EjuSsk9yGSmbK8MJ1FJoECM3Gt2vZcgsL223AVOKKvlAE6XCy8eCpKQqH/VurYE2Xs9aC
+7Lwb325wqqvpVrOoTmi46+KcympMTBSCwSCzrXKMVqb7AAB6mktgOJRQxcA02xMRVjX1ofYwpGI
H2gWVR1ThodDEWvzWTb9+fPYLGQ43Vy/upI5rPZy9EMmNlBQY1LnQgeZFLK0JfP8MKh7a33LhjIw
o+ZbPhHBffNoVEx7Vcc5I9t5CSvySo2/NTkphkEyKt9rupQbMEaSq4xJDVJh1zGc6WpADwdR7WWM
CVwUgAIkGPQEK2b4RPQg959k5E5fS5EXrFJwr1dur/r7KeZn3wRbfYNwTcCN29a0ANrbrJa2jQYd
9I3PT6+wQB5/BH46SIr+ZBBTkqTXHYSzSQLctxTxgo1d6n6ZEKixQDFdloZIPFBIIb3hk75Kk3R1
VD+dWXM35pd9aqKr2dEh1pP9K/uv2V1KISEUZ07YZBBG6TbSSWfCqyfemj1i1N452G8ttBqGitVe
86jnRub3ExExu5eW3k2+yaO1nQ5PTOJZK7ZenQBYF/agoOO63GId5PMGy8nkn5JI4ozoZucIYuPu
jvEep9Ut5hD8m50jwj9y3AxznEekEgAG2pKaDT+Xf0b2ASe+bUWuiMn2mMQpuF53YZ9M/Frhv0y+
NzeSoKvV7Yp2d0YWlw16WEB+mO24BvNgYgB+DqI/zBs3/cDgoHyHqDLhVq0oJJ2FXXt6vXip/wrC
d3Eksy0wsgIzIdoKWMnYG0h7WbZeWbC5wdSForsmkP43Td0FHa/YsGkxGS2SCyTY3kJsAQlNJjgS
yDB0XhJHvaMjnjui5Kw5BO0XoRZ+bxMlZ8d9h3YWL3mQapV/tYWvAnK+6QA+n274Eh2qum/dC3gs
qLHJIRPzVfJlp2TiERQTJM4rvo6VEWyyPxGh4SNl9hr4hDBFwLnGKA99a9HfehaiomjQKEPmuMy1
J4ijtW3ZzguKYzFWMGUQPxScfgSMvAfIPzeNAp8VRcNUAEqrE5bSxO7EzfzXBIcM290kaYciibWE
dPoQQaoP8gwqAqBiqbhGWW436sEnYZEMG8JGi9XqAU7Up7KKDBkcF7pidC39EZjb1Tn/WWfB21nC
tkoQRvGP+M3d6NWxr6i/5lPICyhNGDBhQmcz1uHYSzLQYILSPigKJ6MIyzxMCNieUvT4qq77UyKJ
ZwNi965DjMRs+t5GPaukmsqOglfiwcRKE56w7y4Vc29t6dItfyKj7L5c+0rY/p8IOjmOUx0qbDu3
OOQBfl/lDxEn3h2ERn5HF+++7HfP8h4U8opik+ZP7oTal1tlGAK2uXP5DO/chK5bCBPQdOhKGWyL
HSIzqYhdXbkfwADW2Cnj/T/1VKrr33gBw/tcL5mmUE+3qbGOQ6f9lyns5PLSLh8eRbs1oBC4/LDl
BdlIU6Emmba7EQz2KacHSYP9M3YoT3Zl1KWN8zXGKFkEvdzSLZ3lpU8bYNKeI9bNIz8n4JCKn4nc
mxd8gSQhYeM0MAYc3j4ZblPcstDh2xTrNKUueTI8+f/iNAeVXLp2qHlIwul9CPQyV0y9BTGVT1ua
DCJayJhxZcytRIf07Cf1UHAH6ncNUtIEYTo96uaDzPQ//StuizFEVy9G+z6Ga1v5G5KYgQxxTF46
VXRkPWK2TmgJmg2iWO/dl0RM3WtKALXIQULbT89t279Dl+iY8rJBjjwW1XMbvo9dckRfl1v6+S9X
ds/oe6Z4/I/G469FM6Fhic8y6rf3q0Z/9sLExgngtibrfPW7iS4Gg/UQV9z4fEMDGsBV7TcaC94g
dRbvpYlpyLDb8D6rPIP4qBvrjulTUCIg0YeLtA+8MUUFqAf/MDQkN0BC9Y1XXh3R4OyVm9Z9CjOS
K3Wk1FKAbfT/6BwMcvciTAwxvVt9/HM3vlYWseXEgKoeFospQPcGeGbSWnqY1ab1ezb0bvHLLKAw
Gg36cTpv/W2AHOafgZ4VBnFW+UpQpe1g1y1LorQ2Jfr8gnvXLdGJsAUpReLsBQld69rmc8SU0bdk
Qyp+KK6F+skjeNAMzDtjTFFaLiaA1xM+ZzzmYIHtz4xizGv7dQpRnhaFrFDF5bA68ex+Jv2YNL48
FkwRf0cT/6H4eoAoDe0IDd5YWYA2wosZzZUaQwZRUfESNXGTHsij9DAsyWiE3y3sSjz2y4Q/nrys
FNycxHjVHl7199tx1LqdjNt44JjrdpDFu7Fool8ALSH6F9Unf3vnYR/nUtTgc2beCcJz6j+8+jO0
IBMLJrJS1ew59Ubs1lGh5gyE3a/y8uUU9dxejcwQVdAIiMOIwm1KwrIJF/k5i7UEqeKhK5htfLJv
6sN5axdnzrlYYKnPR/ucQj7L2+m/vaN4evmcYw39TCmOFzfyGDtUGejN0ZYlRMywMVlVEYqnVF8Z
rf4ewTeyuJS67GA7q0Fe5r4fEwfmflPFuw68PxqvtX861+VGm0D69OMaeOndeWx/spNhJ61Ltyla
F3hRgAB40/Ipj3kDxTHh9Ciixqq0PKLPQIz23XOdBIcekoCTIl0DGIrzVLt8/dZqHtsDQrIN/IG5
5izUAeZ5nwdWRRJkt82vlBG7qACUkEZ2jpSZP48ueS6nsykEsZDalzu6tvqflXVVmE3l96jHW4fp
dd9G6jeCwXyaqIx5YPElmjhQPli5XEhraIpqBTxfH9j5FwAFn7SsqlZ61bCxQ2k3in8Hj7WzF4UW
tIqLjQLwb39N+q+p7ysMjLtxm84/29k3jwM+ZeKsccjLZGT1H322AgTZuv0ASiYXIbmFD0nl7MjA
SsdDASmYE9FjiLaBzJMbFxikwqB+IEdJYSJQzjwkHDQpaB0LlGPQn60sevT2LDTUGVZvQwNr2N/k
xDFdIjrQjtAk1W5OH8WFdpcHriQHYXmhILbUiHcV3mNSxg2S59ShbqRC4ZBTn6yZRFoX95s9/ozd
m6orpgDc8xC8xqNw0qFTT5d3bHhzGFkU/GuK+4yJDhjFxxVSS6YSZrLjdXQWPM296SfqfYFg+COr
V6GuKmQhDH2KAxjnphd2ycD6cP+D8r2xuqeI7P/ydXztFtujQhhjPJtdkeR64gRpnXXNaOOYHCt2
2lbHL5GPLdASjV+mn72IOltNRFCeco0kum7wbtOrQtc4VQhd/LXoWbhKjfnVff9AOyyVsrRi9cu5
w+u8r/uhHFQa5xnD7d9/768lcQE9YDbcVYtgejKpAs/fzY7a2bflCUU4eo3bzkY5gHSVlTISCfYM
0FlABwf4ZtexDMIgmv6l2Fu4X+v5qEddQJm0XGET2zOeVcaliOT6ocRDtaa/BW/mXq9H6CxQPbwS
Y8wPoxJxIZRwuxQ6RjM17m0+vDnXPCGEj3LsdUuINCq00kxURU84RiizqSpvv/IDsktwxY0lAX6z
DMKMc3LidMtq4+3jWt4aHThQ88wdrkjg77xWsJyVuOi2YJ/HWnWFO/fqHVMre5LcxgufPqKjxue2
Tv7R0Bt80Hvw5hjx7KjQLwO+0XoL0aNFbMd914vrq/HXwpynsLbbMQ32drKMXH40ajZSvvekJZSr
ZmcK+czcb5iN2Vabjxq6+QPor9RmmFjY4XfF+9c/WYXjSJeBx7A+ZMgzqxg6ezSYg9L4JlF/g2Jg
RHfw5Ef+sCMfR45Wk3Pb3u+pH5QaI5clynrKJ+LUUUMaMHBiNZr76s331/D+bshRaouCeeKdRJRm
b8daDhg5SkYwgXk8CX3XXrlk7UHefonvNaKOCVmWr0+NYHK1oWHuMlYCDTuniCgc7rMazTxIAH4H
/tcMACK8mO7FeGA5lubUCjMzuaAlOLn/Jr/aPW6WMogWVOFLC+7NFcWCKsohq5l2P2tVqKS6LVVm
aeD0RlVaPKbsHse29y8sNGp3nXbwZXjUoo+kre6AUnP8TWt7Kod4JrGkx74r2fYqOl2cpt3z4h1D
15PGJmNyhG+MuaET/r3MfSjiWPYcwy3yG6hii84ATuCyTJ0wwGfAJfMemg1z7q+gYSuXIefCSJmB
8Y7Z5DJzjROUjVEIJE07QqBRY1ORJkVQbLcuU5/KRSbbMHa398EE+xrbfPCuYwnWna0gyc43q+Md
hSXY0c4qeRw8mLOHdbfYKHWste7tLSNXu16sgu4xTsAs6UrKkF5vnb4YhkypsA/OcexwD//FONlq
7/ATcYZXTGdc/zRZQQeOgM+lpD7JtdkrVzju6c8oX1eLMGy1L8gK8V0YxhE67eiFBlJ7mu3YvhLx
6uC0O6eV3J3WjovES8c4SkzsAqZnfwLhIVl0My+efMNG1h1+hjkg/NNXge4jD0HOThq7WUyW5xdV
4xzvyf6M3HbnaRrD/SKGUDpz+dhIKLycAUXo2swEjN1yOGJXVGS9Fw4+cjx98IiFkQpeAoDpgjBC
2d31QNi0hs9o7UWGfaL3pPfE9lGECBQmBCiSr66tiJ0jCi4lFfJEkoYlqJEqFmIxdjncPGzyVxTB
nCzoS17dk90SydgEmNvD0kYpr5SgUuljPdUhR4En+hvfvHWNLB38fgtg8ei4KKczuLbHPdXU9aO1
mzB5EvF0qmoxGuaSdWeFRXhfMnWxRZv1M3FF4NkG8MZhBqrSyjaKwXmArVu1j8KH20bLjg+i1cbS
TvJafhbPtikTlOy0R8Tw8amcVk3n5IDjM25l2ZwTb2ZOkppvIFthnok/MEqpRyAQFX5kqmbVMJzV
x6GOstKAqp9+6UL9kDQB3qM2bulBNPtlck/MMv8mZaTsSvf8H84Sf6pVq+U6UqQ/fMiUW2NIWoTK
6a0ncC1RpV8zxtGPLKm99UpiplQau/FG/NCWbwGrP+kMdNeGAD8UnhvLWHMyTpMD2I9TwmwBA7kp
xo4fS6AKlPu9AwWsQUanWYSDuiho4uFw5SXjOxHLTSAyXvB0FZ4ygTU9irh67ajTwG8YRXQvD2Is
/Lx1V4Kp5zV1BJYa3Y/CIyBDVpqXYJkgfPhrK4glHP4/xiWqnP0HvadKN8v64Ltu+miv6zqvHDPQ
6M4d4WE1/CtUqWf/IHxdCbFbA8Nx2NccL6DrIOf8DV7CW/tPalU68pvY7Hn3KaoJLJZwWTfVL99K
ZgNqR3WPTyrHT+HPQL4JgLv2jxmtopCiBsIEDW3yHP+my1t7IK61dqiGhHR/EiWJk0SUeRjt1haN
FcfDt/fNexyeiRbfte9bE+7EktnaTR5rVPXpf6Qb2tyMh7N8gZ8HHoaTiOrYkEs5ZAhUzqrAPLAZ
SdP/ER68KxSwdxcAZ12N7JWRHvawc9kmCXJXi2H2tcK2f+vnAttd+L3BrP8mCfAdQCOyTmz3GZ6T
55gljnGI8G+OCsC0Y6SYukSAsGieSbsyESSVsPGJt5hfNvQI1liRK8EhOFyFYeFKza6CbslRC6eT
Cosi30TXwOsKDvsGXZJO76+4TSeeCIS0my6V1k7/xShbNI/GLb028YKsBJ6/seJsVUirRgKAOQrL
Ftmo1yqwLmSLNZGMIIT2dTZEZMV4jGcC9CZ93zEdW94ttd0U88hR1CTW/JHETjF1gjgvZadRPRAb
uLP37kNDb1r/RDQ3AcCv7vaXBNgSzgvTX/uDYhLl/ZWMsXDBerfRHClf1Nr218y1O+CKKzGMRgmG
mDfrSyFbUQav/63mN0gjNaKY1M0bULlirntQgrGoBDSwoLQReYCHbw+RWnyuGOrGeFXZpp+sibgF
Dkk/vCwnJLdHVjhDebOtneOGzJLoUs5mKpcXWDcq1La1QZRi1o4vik42VV9Ngs/rwasmrAqG+EAW
7Dars3SH/ePqOMttd/QcbtF8SSyaNtkJWONULsFfqj3pqLuUBxcgNxdSZSk9/s4WGnvJg9kS7cq+
Qb0IaaeNZjyXbDDULaHSlTQdKBIetGBOLRHdjB/7rLHOE2izlDf4Jrocoicf0ARk2ZA+geC2W2wv
jiDnFoidk7b4PJqCa0vcOa4v2bb1cMiT9QsSKYC28U8fEOcEKgxi3pPIezWvl9wPEQPQ438IG8Qd
njXopNRqi1Ty090jIca04YXgs0WUvrtFl3jfByY0/YlwCIB1oD0ERpYueLk8kiq9GaaXlUPwizZE
VzL8cJ35zNaO5xL1hQrUgSJd4nIqc9FAhCmbIJYjj1kNYv8KpRnlMfvABOMFqFc/hta1qbNqsomQ
v9cPYrFj8DLj4ktyX9Xd4HtnvldTaItPbY8swalkAh8VuDzXjNlYML3cBT1+/7MLmuSw0lzLETyB
rCu8GrrzSUPj/S7gh8ysdDyULbS/G5gH22w0jElK8BSX3zO8DB0Sz42MO5HSP7MCD7UB3SGDYJws
Ip7eFErZLKFtV5TCkncfUt5LY2Et/MTpnww4Jq1RVClwxgOFxFz3V2rNJep3LKwCbL9fOgyIJYg9
QMMn5ZZbbqjJ2NVASQ/s21TyY+kq38koYhCOZa3RGChDLxZEf1yYjq7Mx/b72dFuQWesajoeLbo5
VnxFZ7T3OQYANb9MNc4cy/hiJg2p4WuImH+OV9Jur/q2Js66YJbHFcdvN3rsVqzviEiF0Rb9kpW/
4bjMpZpxoojUSxUmkInXvu97I3iRPbAKjTsRAN5EI/aYOf5eMF18MsciCVw1DEY0y7k2h7VpLGD/
5iOh3uphNhPLCOIxd3Dh3dogpl3v42JHMP+zo07UbrgdlrA0Z4o1w9DPlEAUjTNL92a0LJ941tCW
cd3vT7A8aIE3jBpluUh7Jwd2Cl5hq232uqAzm5Ex2Tne7q9UxQ+JTq0rde6Lfcsppkct8NArSgNM
Bhyj7vUoAhjl/0J5yn8Bmkhw3Wy3WVtuhdKyBuNCKqLtVqEtycapfjn0QPIrhIBWKk9VLKJNymj/
Enz8FJuuqV+vWPT4ouKEc/CMgh/MKDvJySexmoxaZjhO/OCo6qDto+Yhdf7J0HpNbO+7CcLdL/a+
h4momxSTq70J0jspGuNcAR4lHZRJsHuojr6rVd9X9tpoAX6sVIWiyHwHp4yR3UJBVfXuLUFfdZC5
3CUSPPcPJattlsO9WbOiPJFyNctngGGvyTiPuqv+16HFgD984kLB3XczbSqXU3d3puESw1W0cZOs
KKTlsKGg3yYiFL+52Fkdj0MX4TgfqOAnlMZ/H5wk7kmxkjILYW8KX8nCFdCEyXSA0uq45lUzVZZk
Vm8p7319IZYLMirWiNgcNYSDbWLhKfN2nflox7S/OOuPFXwbxThroWfD58S7Qi3rv3TcI+cULQU+
zo03wxHwevqFQNMDmd5l/ad7cofiSciBBBQFcuxKRKl7soI9WNcvOr1DxvQgqGoNzB/h8Y6kXTBy
hGpcJ+gEBKyioze5oMhmgaX5S5ecbQF/WaTPRpS66GyM1TYUQrRPjkJY4a5jtWMuoAdDzYm3wIXn
t90zLdtzeCA9XlcSkFFPraMh9YiZ0If1fVmqcDgjh2KA3Kmd+6TPZz/62BKaEbtIzUQXBQlugokr
f3kd0jLibdTkxzjSgBy8NK/Bl0LQXOWgwuuDpFL9/7BQ3QkHuSmDs05oi/VrB8peivCGrjDTsdFf
yAFYKUzKyGOqpD5/+cKTjJI/1nnHkLfml29IEHPXSz97aq1Zg+PY+lZLKvJ29kg+Y9x1psHqzf1x
U/M2RCF/sKPvoRt7/Av/NZQJHFS+SsoMfI7aEbtSWDOH3Y/TWpLOiS84UJXWiEtO6E5qCE/8FQoO
5Xg91DKLDSCSKm+fNCeRNN2D7OC0pDqw6OlhYTrEcLo5dgVeiJOxJDdBoOZ6vmQ5wyt6jdam0z6a
MCFsMeAUxgi0eUh/VQzoQg7Xnxcek1HCB8/xBjB2adpDVNrS4XAyJNsxFH4TA6hO+lG15EckB+Bz
4ZjGCtlahvl5z34z5CkWPtaIUtS/35LVWglEKSsW/7S4BD2GhhpQGF3ayBuQIL23qgGmY6XKbTWn
k5W1ZXGyFYEayVPrZk3GU1um3JOQoL3bI0e0BjYjTudt26WopDbt2y4zrQ8nX9kXB7Jst//XY4Iq
g06+6PTdMJ3xEW9yV5nBqsrcfcboUYwiaWspUZ8EaCKIaGqVI6grWQfGxaxU3IehmZwNc+EBCjsY
7HdNwTx01Y5WxwVwtT0LCENgWBUxnoZQldEJaF3AOUSe+MH5MyvADKjRSpW0ykJYV2hGRSU0CLSU
KKly/CRrUGNkS5/8ZSymaqrFkvKEI91ODcUOtEpFAtSsWtdRkG+k/jdSNtUr3Gel8RO6UW4ihR2D
jvL613uv9C4/mC5sLJmRPj7yNlOmMlaYHQnbvb8B5idz0Az686xB7I8tzUJnj6tx2QLtI6epxXBW
7WW7zEUFPpl5PUwsqsC5Xc1Zy3YnHJp3DYb3su3SfCMpOyR7jMd8zmi4qU9JK+kFE0ZdoRsnEMjJ
gc2EGkLyHN3CN66SXiFl1CVQjWIhKUxMhpfPqZ6071nz8P4AxL2RtjqFOC4hiiuhnxuLz49q+aVB
JCs9y6U3trFXR5Imre1IlQahTeF2V/nFBxer3hi0addIW71WLpZmj6+Jr59YRaFiCD6mhYINsMmT
kF1D4ahQypCfRWPi9kUlZu811E8ZPUfBSF2EqKlOCQXibOLa/BI3t3HUXiyHbVS8JCxGMF+4RjbO
TrhCfEFALh4FVP26CTdeXzbWc3CcCYtdHLYzRmyEt0eYf9yj0Y5WNNo4MRVCJxPGjHkD1/XAv6l6
/fP/YyUvkqX0wx6n7Zhz2pAEWQ36lMUakPilfGN/guHhFRv0I0c/Me+5stSaGLWM1hiAcf6fWEv+
rQIU1gXcsnh3Q/HwGCAwA7xyfBWcadWxsJ5R+GX1A5n4F2fo5uIvATRPuFSUCUNpZ28/aRbuGW3O
eN/Ldh5VG9htDZVTukBWTuMVqPvem0RkVvREm8f/xrrl08KnHEzujOYuw7FbmvofJ5/waw6aY8Vv
BoxBICtXlkBasjKwM7+dMGnletrONZas5JK3CX3kLszrvTnd2a+lJAfK4q6hYjzu0byvgOjqIujW
ZgcXb6TvR7LPigoIRzkrbj+9tu1xP/Y6FjDJzEBDKoOcaKRMkfHRRqUVObIKLAVWsu8en6HpHFEX
oiH58FcPe3/WqhiZLPYnzacTgiwKWe9f0jAtw/i2keNkyGbbj4SV5rif17q2EbEJR8D93/P1jQ7g
1ufZZmBXScKeAcL2nAnsxlMQKGCrHU8K/rALDQ3s3o6N8eL02eqNy83a1+Ok3dxWaeQT2afuXASr
LqQ89ljGGCIICMpS8aT/clThZDhvQP2gpbgraqXIWK1msK7twnJepTqZiR5Aqcj9KBTO6U3aIgq0
0UYvqt0FPKMh05Yf0KmRNlcWAgNMzOYk0qTPQNiUJmxEI632ZSBzEV/sSgZgyWULpyv4WLMB+VvX
DdZWl9eenGFpB6i1LLPw4KezpPQMVBq3co3OAzMRcEJWTVRcgDWb+szAZ953LW4ZiXbSfH3WnPh6
CRcAq0a1C2LNCfTM6YN0E61LJOBaqnTumLDOQg64UfDTHcxeq21Bub5mxYUflqgXUjgXkY8hVYhz
A8zWbkFXbzJhr0LJY2wan/s03mZ8H8DKYafdLL0ukv/053OgkEsXzAoCSzIIQKGQ+m2ITAQNayH5
UvhymJp3zh6V2+SfanQV41JKHUqdVHZTLVt/hA/FUW1UZJvfAIDYmPgYldcogorQu5vR9dfhLf5F
e4DH+pw2hk5I/VIOVAEj8QI8r6N+3GlroUy38cn/LUsyNm2eUgAt7ee1DpTYvm62Qz7fSzaPYgrt
rh0SlQagZa12wqBsMDdP19nEheij2WfOV9RVqHl2sPt0h8hKgqwCXIzlUrcEeT28T65CqrVgnK49
1W/RqJ9N1lfbGXxet88//z+Adpz6dk4XO/XOLYoW7NwD+SjtaJp1QqWiuW4rK34GEnXC45mNkmOh
nyhOXKDcNT+jb1f9ENAq1APc39657PHAcfUJ9pejjA+S2V6WkNi+YvcjvW/PsxHNlbBTRjRTrGGq
+yEeTlVfgRcl67C5TujkaCOa/XLn9D09XmlUphsCvBNFQfGbCBtN52hoy+hZqcVzMgj7eEVHIi6i
WWe8/6X4wizSRFvQeUmIm1B1oAqQ/6tIhddsQNJK3keAsQqyazO+nho/JY0pj+FUAK8BlrV5uWdD
uPk2bgTIz2QgKsvUTjE932P4smYRUqjyOa2jdIskQF+Q6vq9DRb9rOqvZ6tANU//G2rpQqZgAwZQ
yLTHg8zk2vhSOvipWBqmqablU6QEhFT1SzY9Q+oHjkYyclSEG2khB1tD78zgrWeC5yWLLMGrOsij
sRYIS6u5oxC3Dp1eX/derxg3LkWQ/KR2mnBRS/cDdDENVJBv0ANZ4JqVW48ChwE2XhUiLt/mRL64
ZKNr4S3FY3hMwIIjzrG1BOGs9/Lm33Zij7cLtQcqH4yY5Y9tlh2CQgCjvlqujv8nZL5VBT9xpaxR
SBfM8ipciV34+HEIDHKnBF5b0HkFgqghJSEobfWoT9w3DtSWzSxMEpQHf4WaDmrSSTCkyFRxx20S
CcgDqS8yit0QwTIXvghboz+RjK27E9976iOC+4ukeNS9Wd/Kfwd3Ddg5/HctK0+nasQcjUzGEpgm
Zfpu0DJuM4G8mylCkO4hzJGJTeUxUR9HrYYYIHnqaQVlT8m20RaoTyo6kpozsBS7knojkgxH2LTg
70VgxwrVKouwSsFoz+v8ZX8DDBYieBQkQFKhy3PMDouuSrxQutLf2BOeM1K61urH2oqkfJBEiP6O
UmU+GeM+5GgocnTaKOLJfu829qD9+xDNr+SmSw0oikq+GZe8fpJ8Eb2lIHVn6d5xxPtg0db+5xq7
m8s0KlaW3ZfneRWi8CcpEBIMGE0Kah8WEPGV0ypb37R+yhgGLyq3gdXQl+zW/En20/71tfi93AIA
YCQ4u0zNtNZVHzqkbxPOplPiWIbp0/kzUF01Z/2yWTFAMlMCQv9Wx7X1gEpPsG5hHcnRIRYRL75v
2rTX+lcrkHz28J18SYllPYwtD0McPOnaA9mXzQU1OoupEdA/672SCwROpN/88usw4N3xyNm+kc7F
YJd1lPOPLukn644T59pBkKEJA8+9a0R3SF7s9aqy2Kz2bMzKXFP46WJgZbedXri8ivhPHZSkPduT
ongTRmnMu+aqpZ0qW9VI/Gx0GZdLu6L8OEBnRf+231FJg3MtYPkjMACLYZ3uyIwVBfAaLD0s5w9q
8Hepwh/t/LYgZtkipuGySBMLZySE2NYF3Qja+7rLhSEfqPEkin7W65Qx64oc7j0SttWX6f0omLT5
npiSDEHxp7/N6a2ZSnr1yz7D3fW7VWugAFEFeCPFKI2YnobJE3eJec9ZaAck6cOM7s3mWmy63iHi
BCv26Xc4oUA1Y2I81Crjf4YtxmiJ8R8GEswRg9BgjqeMz/Un6iT+HuQ1fZ9RLLb05jHdvXX20TMA
JUj0riULmSVEHWfN75ybQKgIBV9Ebp/G6Pz+Qjvj3mC1U27IBLapsHFgh9U/3Qb7n2W9NuVFYVUU
plOx9VFMbNLMfRi5kMuJN+j49IC8YSCDwpkusEX44izkn5oyfO6StKVZOHlZ6UOLybStCNs7ei9T
LhQPTvRTozQcc0zEm0jRFRPRpTgnKc+5l+V6GxTfbJwdyojPZYCjZhUHysCVKzHaABlPgGPIZ3BI
ydNQTyFG6LwzTLBh6iwqaGpXQ4FPNPi9gr7YthnzQpWqaHQQAFXkKX1j8vGns/214s5oz5U+5tF8
nCbayAKno4RJJDj2kdrSUWXAl+vHM9irPXzCr6jXpwiRFlguooTFCwqVOH3WdqJ4asnvDxrVj+bX
eLhmCW2xob8vPdued7ZxliMx1BD3Rei3591YHI6uYh6RPprcA3JGTIYltuMApb15rVIUK/zHKy/m
jKvi9UZMM4jHqkuetLsWH9TMb2CBbvJuDpZnKiHtBABVOgNUlJCoYyvquqgFUwDf1IrNtFkEj8SH
pQgT9/yq/xrCdTJDmSQhBufJUuKPsyrp59Stt6HP3ZKOQnP6+71JyQfT8FGol2+JxKxGA2Yi013+
aOCTQIKDetXmnbUJv3sRLC5FLP+KasUZyb1rrti24x7HOeys9DKXyHh3EVmagx0wdX8KKG7+mis2
yhqmozGU30UBcWDw26lnyF0Uqe3Oy5Z8LuQueyOfhNfblNHk/Hgzvjjxwo0NoLMLxCOLK8LFfm5B
6rF97FkZb/xiv+G36EVLvsv3UwtVRimzYoMR3O7690ihjLJeZx38m7sc4IXnL6qTTNcDCxbwAje+
HydVcLS0Vm5Et/0vtL6G1eyb9X11c1PC6htqwGoCrIeLVYFJrcSqnlpXv/nGzqIBv6AAEqR1xMfL
OX5xCWogxGnFlFYe6diYA29XSMb0ft9fWloKxIVzhtiR9GOfIx8SWoTtJz5Hx5CUssVlUR7MnnZT
qHri4xEfiVOirrQT3PCDY9xv368dr2QYDTUkiCg5Sxhfa77LFDQbo4kk1ZxJcdQ7eeB164hRFpHn
5k1iNp1KqSYsZX19hRAIMfff1hTnaomUyRMm52Iv5AWG8S0WZmQZDOBnyfVKc8zvcJDAimPh8G7l
tAV6uN687Tts6pp5787Mf9d56VUcXAlxPucSblWbMBpdreIZaaBmRnfJgXbvdoGbgwlXsdNgJbSi
LdAbmB+m5ddB4OMZryrA3ytkOfNTwgmpOLZD7pgCBjczvmLyooKDxwdarBpPG4Fi2IWcRNRD3fSp
tu90At+c+N6OfALCCBWV3afjxgekf5xkqPYOLuKtRDNhR7Dy4JAEIjsBKfLPqjmYY1Y/8nheU55x
xzSxWXMg1YO634heRf6LJnacx4GVDVQjjU7RodWAoFi+W+xt4IF/gQqz79PL3aISpvmnbs1eQ1FN
x5+h89PW9p/Og43vF9rE47K4K159Y04w+vOaEFQLXNyogrNMgxLmF02SrIU4CJAGwkZPtmcXfT/l
PRpxMkJAo/mMQnWkqSnNRiY0JzX3fS8um3K4j0KboJhVhvsH4bEe5r8TOEf6X9DffA4PP4+mejlg
1mpI8hVsNDZEhW+BrtWdtqfEvglba4/8gTVoKfnZln2unGVIpOs4lPQIXWyVX+mjT4Oj+Vg4k7um
fSvlfwbqoOM7oXIXqw/gSNQSm/aJGaXHdC16OeUu/9E8Zlba7HSxZw5FpfVAOL9EIDuGBvN+u50m
W0/PZU9k5zavfxNokg86nJilYNomfmrPsInjIq4w2QVY9mhcgi8jQISXdaXpgl01xSL+Jxq2pufH
6BI+r/FNZ3ExxaUOKlwT+I7JN2azB6Icm00zRFOmnQ96KrQnw2dBAiruxum7SMjAholBe4Bh1gB0
uIZLI6j7ywubdFBaOxKDJoAxvUzI39xZ3eZx470qncJZIvYaPabpzkLYiDoS4zPvMPxfRuUQJd4B
xLE+q4Q/oJY9PbIhllngDkQOvz1bs3a06FJFbbK3E0QA63IErMuVhUPvB+qa2PaeuCZ1pW8FWFnA
KYX0flzOb/bEeaBl9os7I7oS+GCUl1inkiFeVRMaKvE5ujyiWZPPnzV8+XHSppu8OE52Hl9+aQG3
zcaoTgJ85m+hPxlYEEH7sLtKYhNJJRVsW4486SppezBuBkheOaLpgnUeRtoDRUYR2r56PmgCeCyx
QMqItll33pvY/KI9Qwbj94icYzsd/4T9WXJX50r9PzDXTt0sqQvkJbIdvO9itfKg4ppvTaGOMgLX
jDviFIolQ4lrBYnZuu1R7LFlEHcK343fofUUd+ATzq3IbEUIwW/096gT01g7YAfxqIfUa83n6Bac
ZG1yDDmTuPWwpr6myX2QGhbGGP7pzYxSwUgeXtqAPuv89Jhx7sb+T54yDhrgO+dej1yvDsadm79M
VTIOwjK/IfKZCIfo9mV4QuzkBHOjjUHyXUFX2qCIJw1w73aZjtFQ4SltFHJPr2zc5NAClpHfQiKr
L0OjFM4937IOEGJXKqEFo18O9E1VaTrdiI4CKdLCj8DCStudIu3O9PQZOxdB1fuhXvlNP1EZTRs3
njtcKfvglyOEyw7ykKg4sLz6Oxj3QO7jl6JomC2IXQ+o3mb4CP8soKk9MhTBOz5sukDAS/iiyRV/
nWmR3UxuBxGA0dYgwgz6chHFkZK7PidhYnsV3uOeHzq5NhBp+oheha2W4LQoKuO6QkowDvUY24Cc
IQ3jzEQsjsIbHN8esq/y64K8dniiLnAoEgEVkq56Lt3QY/jLKmC0uUEkpG/feUe+1jhoWirlKpTN
kGAO2kWSouUGodqGHEo0hx09Fl9+1bmIkJ8OfzZCHH6PDH6b7N6t0jzLP2QD1a/m9jhed7PzMw2Z
wjm65+gMfxlg1jv7apjHuurWNbIcIn/T/1Su1GK3bGNNXvZBCp8CQWOBC1VaySfCyqtnob2dRCR1
iVmKPs/W1+QndmnRMA6/gnxPRRu4/Lqorutl6E2lVTVFFutXaGUJfTuI/0OCi7sAMhWd2arvkpcu
QRbbwiyD50avHiFsL4OQW8yTa4yB93VbrNIhGO/uzPlHJYeuG6XIvx4gv/wUmcmbDB43RqShKvvT
7PRjLcm6JELT3TuEDop2LsgLy6eDOXAxU7YsSZiVt2mGUYoz4Kpqzq1+vaVv4ogP4mZwZHgRs2G/
Es3pwvYHChrNkjAaW3K7LgkeXRPl7rguPrOyPBid4f3YpHbYiinenH5hVz1Yo2n+jdfn/b2xqdrq
KmQQHKWJdtQU94nVbLd66nc+IFz1RwfgG/gJk+0x2L6TwzbmgyI+qO3+D4kkUizumg5ZHDgobvhI
ByayogP/SqcZ4jI38uIxFVkgDLkruNuh8jHp5xbkY5oQGACtA97//ETBlGW8rivikFlYDBNil0hW
h/vH8hJAgOKKz4xhYRafpomhqdrCfS72s5yTUaLkI3V93HtMHthlxpWZweBnL4HEUSMWxSCYssZ/
xTraWi+97QOhJB61YRsSksVRj7vn3p6lgZwEaK2Gs36F8NKVIQrGKS27mXIecrUXhtdWqJziCmjh
sxHDBXRGYwRsQB82mSNcMfDlMo3xo0Hs+VmVz12C7o4ZD5EKVkmV7XGAhPJdy1DHKFEyPWks5q72
dIaxEWAZLGhsvTHkbkI4WGnIJ+zR6nGoc3r+pmb/pVhqhpom7W5sWAuxVoEF2aDDxyJhm6J0Xd5q
++m3xzCbpfbpoqjncXVCrUilze7QTnZL9TRi5x7zJB/6743ccH0oiE3YY8jXZJqZ7FIPJo30RWJq
hkKOFGB0WAHFvxj2lY6kseGzajvuL5o7u/V8imdY1OmDuzlqB5wzEej7YNbennbLaC3BxzhB2b4C
/nnCu/XUQYM5y64vHTCrQINJkKeQAmvnPyDtstlmVTIl/gnR/VY10KdFbnP8jFvtJbj7PSjxwAaB
Tg4WNZCbjBmJbsc+DpyD0ZUWGMJn7iJ6mbkYUz7cokpFr39WokhWDHoQBUzp0iWiPdcYd+GBw6JB
V5bqhkYKsx5iylzASaUjsz+q+MLuYeBFaFTXo5hgHFZOuH2TlAKw3QRpi2F0c9i3CUmO4K5NmZC1
8B6cozUdZFVR8050jpIRaDX013wvLYjvsRsY9pP2v9zgyNeUZEt38asGBfhIwU1jPFEixv47gMbr
BSx804nNa8V0st4vm8G7ibEIqIz6pLzHfh5BziHURt4C7mxZpJiWiIO/s04kGwGAnijIF2lmpS9E
96YsOew6X5rQOAzla7i27NRZXfZj4fQ3eosZ8R8k0Ryn+vMvi6GY4CDQaEQagtmDKMWKK7SEJN6n
ArD2+h1DnVKKplHQnyRuXeQdYFSgn7W2FkY/2dFRU/9zcgWBVOxK84UdWLd0OjSQMVBuHCcNfr6x
2r8XuulrLvSZgbvDmthlgb7jWrBspLlko4PaWaOMNEP73N8aj2bu9do8kBHuOcpd99EgNSQlq8Mh
5lo/VmbfUw84jP0yYcxIAkb9q3ElZ3sQxwVg8rRQV0X3tBWt1Jcm31MGn1XkidwE8GZRhWrwmRWC
DXaurt8VhTYpmaIWHyi0Oo0v5T3hCqnI5/mLaVpxPed08qMkym5HY66NC/kBB2iciZoEexr+Ia1D
3V77XGgIIj6bSBgH+VHuanNdZZVtIY9LXRgNMd5WBee0DQaGLu4X0FKO/J7g2dOu5WoI5cWAdk77
aZ0J8m4OuUb7OU3X5vP8CQIFFZ1SNN6YTV+jfU6qo3nIwcX3HXzFg/suPguYdj00mhhSA5xlVpFV
hdLwKOkaHnOhTuDo1WI/msKqDzPsYoGeXH/eUw9ELOWEqMMuVGO0zbDDKxGpzTXvEnw20Hqe8frm
jEI/V1uxuwPv3Dfj5RqFbK8pVwt6Yf4mPdar5g15YSE3fDGKI+9Lv3fdRekrIHK9mjJzi1c3ps/d
WsS4sIEQSwKGHHLG3n3aHCKY+A9hnEDFz/HBNUPeuxm9M4vskS8XDYFLMpo5SQoTfAs1g1FVDqOZ
xQ2F2tApNsGr0WDhBiuQVglAQvlZJXjIiqONxtN4cA9ZVW91THgPusUO7w7b2fDd+MEJ7SHZ11YU
uDH3o4fAEOT+4ibXvi7FVYmjc2YezcEv3mgvKK+GieIhg2h/BkxHFk2GJ8DWjFufQ8Koeyny6jhA
DCZs5CHKVnUH4Bo4Uf+DXD8miMmo2MFPC3f7WvS7+UXsdhN4hj2PpxAx6rnRC4jHwyqeWuHrPkda
EgCXYUdWv6XCyYGlg3aiCIfhU1PnpXjIlkv5TRrtyvtqOLgD4f8azNI8NiC5/lEIccz4fkTtiBPl
e3VdmkZA9L4wt2L+zk0UZm4nBcnLcZyTgRYE0qADwqvVnwTJRROOHvEsVJOxtjq9hF1mT6isPGKA
vk6JTK3tVX6jsvYH370JTqwyHpgp/K/d8yXbbh0UGras2u534M+y5CEBHmP4x3IK7PnTT0YEqsGa
SmlOB58vZgH3KrYJjgCvQZe2QTElOK4642J7+YvjZEIgNQex8au0ZW+huXhqR547sZcIxC6BglUa
8unfEwjaP+n0qi9/wxK98W6WiTaDi5Er9/03DaYJx9mrhIIKW3GCUKfFTVLhzbm/CDlSZ/EZ/NX4
U979uLryblix8pgc4haz9d1WSTaxRWWC3sqqbDmPbsgtfJss9Pl9tTr9wepWecjGJIeOrlNQ2xtq
h9zVZi6mJOyALvz3GjH1iNxkz07uB5+1FEsiJtl5dhy45zfnX61GQQ9HN8Yg/9CfgUo2c1rSVglL
MZo0QNzvhw0RlxGzOh1ViTUgcL0Y4h/S2/xzvgv1WRPtdVyYXERhvhQt5Fh7ZY+OgMASUJ/GbDAT
P+HtI3NwF2wjZjwPYKqRwDqq0RwK0Y9ieDWcmWyY1mwCNBB4OVWsc8WsU8mp+Wwtd8/AItDk5cRF
ZlsrPHjs2OOnqdlv/eRD9lBUr7Jj+liXznp5fJAL3bXEOElbfE/df0OnxIZk7JJuQFn/jZhL7MCm
xMNCrqvenNkNjBgFysOdEPAGre2LYmJkH/VyDbuH4kyo7AkWZPoQ3hQaVa2yW1D87vzChO/Npi9Y
sZlag+br39wgFDWbfJrL+ygL0WqJkfaUwhGL5OOrDhAH/NGHnh0Li8+aqnlXFQ46JGwTWIDM6kDm
IgR6ZUNAuhIqM9e4/2D1XAp5g18aboPMofsX+WGy6WLFFcLMAGEU0Q7ZJGQ2Rqqn7Iv+XuykVDNF
1jdoCHOBVqDlHk7AxoKqlsRC29sB8ZVlNMUV7YV0EhXQk2kM/IWQVFzSf2upqCMcShGJQe4Nq6aW
Jvvi1DqdpfA8nK2i5CN7spcMr06jUE7wqRBRtIomyYMnYHYaduvp37YVwx5ejfFSdrRPUw0m68vi
78U3uWvsA6/ctGMQxwX67LDylMfzIIG7LEOb/xFNIDVXgCap29GPWOfFJzSdLyyAB4CUr0R3ry8v
lxVtmp6UpIuF+H147OLpjcQeuD3vR39/E+4CH3zMr1zEgSHoMX+QrR5y90gAxlRWhryhS1FTcDMn
uJlyqyrV9/BncNa/fXIfTQ3IGw9zYFbD4LJVfmrxoX1DjcO0lyW8VtXWbHNWqUI/tJqLwM5ZM1OR
8VW6lT6IryAsl0vVhgc3lZOk2jcBPlK2uKpc7YL4yvSxi3mKPQEKY3NVq2TWkJ41McKKajt1twuV
HRxka3BYPqyIQlOetZnbeafRgTyCvGHqQuJfwgk0qWPW+QKzDJoOYFrYvUiiXW6D9+L2E/i5D2eN
pB/bY3xZjUPCFW3ZbsDoq4jxIDTdb9b4zEH1aiD25xSkU8ZD6Fl3Aansuud4cRDPrqtU3O8ZY2jV
Q3OjyEJhPn8mFKPYrfRGOTJbd/zt60jGViUaX2ra0K162tU2BhOBv1GivUbxBd2wB7UDqb/V1Dht
cwtGu+XF4xUz5FCqteMGYzaPD4+N/7+k5I/ZLzWOFQP6zXmak93+tjst6DXkfQaHvKjGYeUKEm+2
2jI2s3fkcGVfNghxc7neKQ8/5JFPoyzdeUehgOrHZKHhdcrC0aHHSG3XM4n+A38NcdZV6paohXIu
w+Krxjg7soL3rykhPwYe6Jg5JCuHURTnL++r74ras+qxkAgaDkdLCFDApon77el8QINpFDtxvqyh
HFWK7qloQJG/UyXiS9aDud1Y0vZYYhBfRqUgFWufQ4dNzb4qiY2dj+jzpPThb9yg5d0xMFusSOQF
viGVKUp7EyCM8m9rCBzps/vSOsWb7T88n71nMxy8HMjIoyMiMCHtbgXlYSuSR0m39LFgfO/0izS2
kyIhHpmSYROY+3H6KRkN8AyCOj4GBUJ/IeN7P4qRUlwl/LSDhHC3/nTwxnIaAhlTzuhCSJuFbW11
cyu1MDWaXnyNpXJ5XvnqI6ZptBc9ANB/219v2LPTmz30uBF54eSZLoWdNpHL1xcOpJvXyfZSEcie
tgEMQgTpSTMqVpHaGkXGUxzo4bU6HAYZp69MUCT5zNO6bwgGW+3eTxyQh4HQl3pT5azDl3CAq0n3
EKDsF4eQEeu1OnI+o2v7caaqyR4E5Ek9UbEntuwrYsuKAH/xtI8zOUKyfRxBSenM2xQZg/ndfiI+
xSo2q6u5PmApr/PtkK3GPXuITuM3PhJDWLmzZjJ7zovIFvLpeY8/AJAeS+HvFTGDFMqGQno0c+1P
gBFL1qNBFbTxKp11bc8j/hDUvLapAWx4F/J3h0NVczZar9C6fDypO1WY8T31sSLZDfamiyEcK4bY
7bTocdmzetf5PCxYpW1aBJt9Km0iZauUpZugLTu6TWFEYrZ/9c05Ui4K/nE2Jng5nLoW6IOp6Fv8
Ba96tIKAfGNN7iqCxIalejRUjgDKNvk8/0FN+tvaPEBwGBcFvlQjPJZW8RJBfIYd5h/+0vSf/sod
/nJVWU2vyksUvq5M8Rk02s4/VLz8J93/cMK5YA8t/PAJQ2iu4PrHYfjTlEY+zlTe8rWYvdCY1BMA
oMlUEqGJ0A4GdN4+yqXI4+sG9zM6T7YAWY1gtPyP3FH/SaAslh9LIIGnQiiumbFvrz4Kg3xXVAgk
6OzJhtiXygltYT51QVEIaJfFkZkqaeUqmreAP9aK7XvByMWMZZc+wlOXKFZ9F7RS3Aalsv2VeDNQ
Z+BAyv3xdcqGbDU8NBAiyJT7vMuN6slTOZk9UJfiP7X88bGW0PYxpjh1oz1svw0GKZ6XL5QBuCYK
TCI4gTAttlrpiHf4OuImsUP/g35SnE96aFWIosYbmoY1KkffT8XDZKLbduIGtiE5/+3txDeuY4iu
ZIURXkM8cD5RiCGG89Qzuwn3hR3xHsv685FjEEuPgftlRLjayiC0kBJzaD/HmdIxFRZQIWuJ1Ky3
D6oKyRRgBLSYfNVj9I7fOKLKsPzchBI1ZzM5BAYsrrcStFILHq7d8+0ksGfD1P+Qd9u9UPnJ4gVq
ExGRwCvQr8WwmscWMkZ1yv9eck/RrMiTbOcxs5T4MfQIa2xqI+KOrXARq1GhBMdCtqgi43qdarPt
IpsyPI105S2kUII6DOmpXWqZrGXwIBX8E7ZityBls26hN8dhUVeAyuZt3VXFuJutMS29q2/2gp2y
R9ueDfGe8wapkfoMZrpXEZ9zyLSc8LJRAkxw0stbgI0UkauvTR6M9ILGS2eo9OD4nQuUWyxV1rpv
yBmLfYn82trQ+gCqYAe84PXBVaNw4l86KFNTK5fvqlT3LNlyYUI8AQYx8KT6OLzBnAvkAbqTbqe4
m7mVzryVI7INnJVfidBgHZZy6Zr+f72eWHmYYnhepU8ewyq7hG5nJrR8BRPXyaM249oVAeQzGdr0
4nA7dhaQ0CkrCLwmAn2NPC3CraOfrhvxJbIlry7oY52SQOHx7c4hsqBBvbovIVWMUXm7TE7VrGna
eNmaBTDRCsVbPaAdoX60+96EmhpEYSMXTSkdnAEeWObDAq895sdwFHsBK8g8b1E+8L4k6PLSHkPs
81KKvZNkYEDCu9KDm8mEWUR0po/Eooetg0tpGdp8wc+lGc3BC7kFP5C9lC/PcWa6/VWb0HoguODm
iqrcSCR2rwQXCKNFoAzf0POJdZdWXWzUlIdXJoXWJm+z4EIcyeB+r8+5uDUUcTLTdPIB200JBFJj
1aElLXNVPD24z5CvvLZ+OMIbByakgxKXxEtjtKz7QUkx65WWtuk+9fV3+wb+BAUltnTNQZUfRXMm
wE4fk88kjYf/qQeGP8rjj6hbJp71ZvyRhcNphOVbMfy8z+llkFr7XCMEbdBosakBNlODlhIZqXm0
ZqZINVfZO/DUnO60b+SFbZb+XGI6uJ4ckg++ae8mcK3MIrUXVULP+2m8CaZP2C/9GxZILapIiGMF
hTyqy5YbugZYLM/pzwx1osVa84D8YuLY6AYUkNTcJzIU8NxUJYUDHl3dMeN4kNdJenHhF8+nynp3
+mr4H4fT8uvHGmGzz4aIQSHofNio1wptx5i5Wvvxkg8VpNaMZwLjlKHwywq2QoPbW/TUkT8I4HNZ
o28Dbi4wOYSOGVNwIejud2QAgUhzsNz9zluGuz66Z4AVspBQxwPX1e+5BUp4RrTXwOe1dyT09vSH
AMmY0oPNzc8p5urzat6Val3BrVzobb4l/ilYE186D4CP1MFKb5qhI1WF0HN+gT8UYOpo9YiRtwoe
5nYiCIvJIgeD3PWIvwukRf3SANmwMN7HHCRBpLlBnsOdIsSLb+DpUektZWqAgK8Jds3/8bhQz+cA
ELwWTj95aob/5R6Dz9hHLhsDI2cvWYIfRO8s57rVSAPGIyCIEn779uCeNOl6BHVqd45j0wWn68tw
Zgrmvk50mJPZSN6kwDD7UkPzJqsgVzKZ/uapR+JcZY7GpQW68UbqzS6ZTgFTQ6BLn3PSLCLNGvNT
Od/qMf3efSnNJkFvaRYOtCgeL+PjMuV4MCOOK+Nz6f38GDGuMwBE1Dhj1MLB413zDnZfxXjxFShe
y84SSO/8IQcRb/1MRf0aTNOuRO76JdmC7HmGYzWt3VqKwLoVRkVfJGzUoaWaUBhETBzjvgIEJiAS
vP1Qpikly1wcE3Qx3okYKh0gghECFYQHaYdEzBiPwNJ0DN9GC7eqcmVj2r5PNgJVcirfhcJwhaiy
7lASK63ULbmXeBJzQycHepoLtR90VA9Qc72X+GTU9S0bzgAB7URLjcf++0gxrCHCwEIQrKIIZtNW
727iFdsT7sueIcgjVJBISE3rFxB0IgKnlaHUJC+IEcFq4gED0Tjk+rGpgHnyy70w4mgn2xMlgm2k
dwT24d7uZHQuGQd/Wq4jJO9AfKwtY/A07hN7neMXqcXc8eo4okLl2izRPb43qWdHR/X150Jqk9n5
49m/rqpvs6Ze82qumiUSCWdx7noNX29FOt9/A6QZ6d0efwnNqykg2WMW2MD3s/YadSQ+j3Gg3z8C
Kz4GBsQ1mvmVoUECkPMyiX+Lcdzcc5O59/nPzcT7WdKjyJA0rD+CjBymEoJscCgrrApMVJaqHjOT
5eYzgHhAdUjbrxaU7/gx3QIbJjYGtoLswveMNVJj7LBQXLofHjPMBCOERBZAHYPuGe2YLas5Onos
Ek1Kb135OhX8LDOq78oEwrSLHVTnJcJ/utJGRFYkcBSWIsFDS3w0e7jM/5AZyXB7Ar6Vc7lGruNr
PXV+zM1tiWc4vHW0KvdPfRsDIyOXeE9x2ecqu7tbRctuCzQUpOBYwvR5xzAoP51dnYI3W2cBBSdU
Iv9TQ2220l9iDRnn6Ni+O3iIlikaxglwJ8/ocIwLeHNnMT3FQhTqYfvo1PvR7jhX44xzAHa+SYve
SPzurAMON2nQpWKXZjt194/fgpU2g58RNw5cx6lCRvezCZtYCdfgUwALe+NEMaedPtQU7Bia/Jwq
UZ3T+eY5xMMAk2AHGDa1EccgxAGlEaOqxsQrzLfkmRkqJA6NdiivEvSlfnOgyLMv92sis3IIRqQD
lRUrPmORygsKsq4zS+k8ryi27kTOcwIi17i0XnPwLPre+Q78S120ibqoNyJgbxjwpk2A5raYeUyr
fCq1QX4fOxltMgRVn1Hi+ixPzIP22LeKxMm/BQiEMrRzbjYI9bw7w/xTiAZ2ZQQ2vIXltRigfmX1
z28spvOjAhrRMvmPtikAIoWxCNFm3FLowo/SmxemMe31WwOHBtMJYAr75VBAqqzdhHqysvywUOAm
znra7R88Si5F+kgZcCt/SoHiIfqkE7xzwt/akFBzOD7dLAgEX2mJM8Y9nfXdwPW9YH3lm7DvUQPM
3vD9BW35ftbEQ0FMASFZ/Rij5tNT3i1cbaCUfdbC9NMw9Dc8Vmfa2XDUpMHcaG2eLUXAjKNfcNgf
vtpTN9UeSM5sjOP09vKD0C994/WC9Mqlddf+mgr7bavfu2VuOfxyt6ecwjSZkKefQTXOikvFxRSX
QO+wiJFJwMDY+HJM2Fho5TFsKL0ht2WRqL9hBhufE6yHkNxU4NSz+FANokDU5WgofLAEQvHUIc59
I/fYV3Hyczzf11oE2FcW4isieVCvTqcwdhFhh0hSKdmfhKO7H5bxK+5oJAiFHycvBAomSutqok+7
8KJeKrNJGl/rRlFgDjoSBTNoe5etlPgO1lls89nj6T7z7yJDJg8ki7L7tQkZ+l/M5Oixx7vAkf6V
PrJXS44bZFH/UJcbt1OtSmokhYOqu10To+yzzdi5ywWHYkKjuZleXd2C3y5xyLBNQIV0D2o+bko9
jAjNn9vCi0ZsN1V1pBYoGAw+cvBtT66ELkRof+vQEHX1LbvRQdn5GuZEQvFKlJRESjtlzLwEKR+K
+2YG2OsYtlK92KaKW2YpNEjqhMkI6AQ0BSissCFBLtp9JFdOaRmnnQHSD7MujQtSA0N6WmPQ/AHr
VvlFwvP4vAK+yuCbkDi61qxEqncIvUBdyi1vADudzkmE5fSNQwIby1padRr/RY7t0OV/kP/RXUSA
+QkaQqW9W12m4Lsl6bAQLsQLQuriZ2IE06IJHBp4Nvtx5wSHTaZM/QrDMPX1YbHHe0aFVtelw86a
89PDMCXQfCu5XaCTnEeB7gl/DB39CjvFytSvdBiWKUh0SrkZLpfZU5XH3kvaDm65AN8hxtra//NL
/XitMhUqN/xNQcyAhrpPOFqPbPxcAjyhBb9LgbsJ1EABbnSE0qnPSbf7WD343rB+IeUgiFGKczJW
Y9eQLDv/EAtcvwCqqm+o0aLB9OccyTD/iLrEVgJOYtl551V8BCZU7F7gdSXdA0W12jgD15II90sx
yUeJwO2Ii366tVhy9vZfacgGlV/qb48Q1QxGgtfOVpeh7dUIrAggmW0Cuwe+aNkjDkF91npNTn59
LjBafmMm66m7wLHUCCN5lKPNKXaiWvInBCsfxoz0mL7IWUHyJ1auRjwUTel3EYLwZdzWuv+ATeYA
Qa5g+3I6ydbmW+buzta8DjXcYf96ZPQBeaE2tXTROk6RFfp1xvQg6OHnTseym5cLgFtamYpTZuMa
YMXWlu3ezgSCfj8eHv1NJe7UtpvSe3/lNudpHEDgRaSN1wz/c70MNGvE97pdDszH/C1bjiH9H/mf
bZzulDs8OIl+0koN2RFcXc8CubZQC75Goc+09btaEon46DPZIPSNXoBNibB/jrSqU77l8y0e5+p+
die0gi1jnIuHfZZ3g5UvGM2NMQp1KBxr7x9s4vziKZ2+IFbM46iAF8OjiVINmqdkjUjzNX3DHxCf
PVP/SqwTHWPCcdFDlU4uLw8o83W2wfm7OQcmojLxLDiFqr4Jgh63//f0tXAgbMY+QYMt2sM8WVuS
rFcgNfEqZtxUJ9SQ+abT5BtuCMH6jbJ/lnRUap44epTcJNKuj69qONfHqUq9+ePhuysEfmikb7Jj
mIlc2AF7dJOesqlKuY+FZ3f5LsDfZoIxTVhIcUZEn0Onh3ZirL0Z/iYP6iCjxlZCttxeGOON22/y
LyI+8cgiNIBJ1qdl+hNE1ZIdubDbKjNQXWsc1b98Rw+JLv86glawaxnTgFtMuisCRNNA4orrtQnI
ZcjwhuJv0/Hr941DtydYuiNw211kp3CmrLCTEMvriJPXUpTlVjuEYzuln6WmI52Y/VrWVPpTU8Ta
C600MKXK3bXJwTQFE1kmq1mkdisT6Vzk74HjMSsL60RBTPbpjZzpK+SWOmtF08NqYQgXoS2kQXBf
TPrlEfFCzP1dPKVDdiZt562oKKMxJ45CMEbaLhSWScJHEOX3KhoBc4Z1k70ctKLsRSIblNqaamVz
HVMqMgwE48N8UPKYWKBMQH94cgUgye7szE1IDER1mHsG6gLGDKFv4C7vht149jxeWma5xNeWAHJA
KdPmzYhurF8Ce6eOP3NRfXhPnGqCXEqVK6ZFNDmU1B/o9rAbftVTDQtvwr6sBARTiH9knum8kc+P
HSoDKjHbpucZqzUtp1NQ+KjDhaQMHtqTkWNcD42SRfye9YNarvKl1WGqfKI8l7yRKcl1sbh/5M3k
NbsejZcfv+KVq1TLKPHuyXZIoRvSWRi4EUbQ0m/8yYhpybsGPCbY4Xwu5rpxoaAksvZXyqNVIcxf
tXqoyHolf753A3zUi1JzzITqSHDtJS43qIN2t7qf8CA37frX3by3RdGoqkZp0yz5/bO6YNDNMhQE
XdGVuFLm1MkRkgNUeDYyzEBUsYMHSOrAEm/flzc40BaAr4pY9c7x2ckJi8jIUFZq3oP/kjAhhgBq
ENkQabVF4aSb11Dinsepi0QTTtEiyxgaLWYsngi2k5n7/fxPfQWjZVnOo7fcSL/74Bxd+5GF+amL
R4kXs5dRu49TflKJ5nYKR88/x5Dr61CzP5aRqoX/Q+x2zFaHbThpXagf0/nBywyTUauirf+uzeHJ
zxddsOs4J8yn4UHeEwDcKDdI1bTbaUdYL/y5laTEleYDSUpKtXNEXPhj4Iven0D5RY+Wli9vaJ93
8TAVO3fYyO4gaxSw6OHAXV+BH55GnVGPlU005okAvahbvTPbL8sDRZo+LpoBBWDVicAsC0vxLGTC
W6buHOjGeEfCDH+mx2CSD1mA+bZPi+liGYQVG2iqFjkwybiTNaO6pbKc/tQJsSKHh4p6rHXBd93Q
uiiBDCzeE38P2TY9Glgh82jZ5vOvxDx4GSA05WBh8RZEGarO71cYbyIhYHmfdkAHS2PD+7JoZ8rL
WQ2/yHXsetvQQKQ9GSK+FY6kKVE4/hLPYvaf9QybHnuFcIKEkKhBda7nwHlWUjf7rbXySxgVwr7/
GRR3TaO0cdrG0ptMhykkH9SPNELDxpgLffcjk4c5MVOUTMvbNfDFk9UsGPy+hEuzo2rK1WFwA/PX
h8f/9iiPaYmC6RCo6Fg0T7AIoaBrlNs5uVNq54faI9HKQhDlh/TFZZ8ilNMaUszNevK6GhpWhoRz
hB/+4aps3q/1kg6EqAbvUtVEBKwReYY/82jlGrJRZUN8osSdcYa8rnt8BhfIZ4twFCt0OS+iaNLq
RDvGDuAT6WYZkrZCCpM/ht5rOOCxJSrrQ+t7wHPJpGOAoZrMI7QHxY716P1jtKHJ663wq4xzHe7u
oW0DoygFSF7CBimTdmMhVtgr5fz5xC1YmE+yanYhHRqcOGdPaQuOQbY4RUhjbsX6xAizDIptN2Cp
/SsREQCS3nWpMF3bxLlzSV01TZaUREbNselLsRKmHYWC1+fqhoBzKm25yPJfhtcklJn5m8h2v8Xy
dHQufGMsX5uSDj/OhnImb3YwaD7B8jbA3eugOm7QNu6Sk2BNbeux3hWO751xsoli/1eQhTdnm9HC
wXZNOnMow3etLKTzfxmNX+ovzi+jiQlr5/dEy8m5L7as1SM4awzNXkuuTesZSoKcVl1YG976qiCu
Nd/r85suGP7F50ZQwq6ZC1a5oTyjVUBvNeWQC4gUQJ0sxv1rzIlzL7ywh7QOSpQtx7V9J/g7mMel
zUiBcNKn/6PQcLO8UFs4Di805mEeFWGxO01AmMsr+bV/oOk/2nPdsnrAJJpIF4zGs/3q77pwtn2r
96yrh3BZ9W4nNGqyDIpXU3JnM1+nEGUfWSRCcP51SqDod9VQ0R421s8+dYOF/7Zb8b164/whxUGZ
RqVTSnC6Ysi+6+8OwjN0buRo7e4efyIJKB1CfqFHYl7DeHHW2HIPptFiqCeZuYWvwJ1WtGP6XLH4
gwK86W6fQftf7ZTKaKnl6AnEDqToxlkOFejLXI25ykVgede1YgFPEgAMzSpAurEGRCZdHjeI02+5
tncGRHlS5yR+8WRhcvqETCemMdc9ZcIKijbG/2t9f15sc01ic4v1gGwzL8mEMNsJraSRh11+9ZM+
uH1CXg997Sw/DTBZ4DNle3+TF5EHYhU/4a/hBVy/4Y6jyWHzdhXvtcUklx+M8e80YVzmoEKsuB/B
zBrKXUL0EIvdWqVFaChk/9/UC9ybG7btGFXuJbbOLKblkT+QGcotfLm92RW8arntAms3v7q/nXl1
lzwOrDJNIdeMdFsVwiFjwyhYKSROP2ToFPwZ8hA0eCwqQC3N/xx9woLgJYHhXvOPIkqtnrxDjLHd
ssa2kYWbCA7QpHyqvwQcZ8tM7wiLY0FUQoQwBBFrWRrBpL7dwB3Uqx9H36wXLBok2anps6fcnojO
1VqNLYo5bTc2X8kIMBw0SCdp1FR8aqDTtvX/VTnANL2M1VNBzGEz9hJ2RnJg5iYwNqswUaY/U3gx
bju4sGkzYHnMZeXvz2k/fH1/eIZGwA4dxPuAceSQoQpBETm94Fp1WGf1De/tlqJMRe2rmJPHEd/s
OX8V1xMi3Oawc1cmNGTJfCBw+V0NOXfgzCYcXnTVCZxgoQ4oyRgopY7bMiayVqvpVv5j24+Yn075
ThE1iZ0gsuUl9QU3oxdnk38mXC3WlDqg78NCJZPxtX2unpYrepDJbtKhtyJLMnh7PxK0Y0pWvQsx
fH7U/upDlyYZEscttf3fG1e8uckjQLqsZQJUD/PV+Q/1IthQ52kxbBoR0p7WZnC30T6ZXuOGPZHx
HVr61IOgHcqGR98B37bLFMlxYlQJEEytyVZDaAxcBhLDkz3P0VRbz6AiWCu0cRMjcoF3ehNUcmfq
yC18vPzUE9XYkkDPuQodaaRtVJW1++0yXQF5CtgJbgLRjuckS3fMfK6fKpMyr3P6Dzt12T19EZ09
KBYUdves+RrcfEPZ19RpQqc+t3ziQfQO+SJMJK7ID4y0LdPCcBt0y3ZBXxoLCiYycWMPYx440GK6
PGmVwTNbOiXc4/32e2av1ijPQsy89ms4Lss3bWciILtewKKPBT05w29uDb10J2hZtj/rUcl0/V7c
KeqEWKfB1kRzeP+3fdiGrp880JFp4ITcCBDuz049RjM5hB6NlxZvCF9BuIB/ARHnk3Bx5MNFsYLc
tgwYyYXoUfT64DlU0fvZ6VMJOyfwIG0NFsDI/7RA+/rHOprdZup7F1mZKzdo+TTfXcV0wI9r0Lj8
Yp7P6zgQyQ89FjohGqFDyl314GI1XS7f4Lgdt2kKWpGdFg2hfpv6aXEUrLZdECUrz7Jxh2WD+VuJ
/GW/1sqcg22HWUHAGsxRGXN/XiprMgJA1vcy3s3mp14bZjJ6ar7hBjZdkdVjlf58coix+9PQMk+/
FXeXIiyLuYK7cZXhujBjstjTJdUNdUKyu9JiKt6Mlr3juKn0TPRPclriyTszzxIi1uoYzuXpZ2+J
skxUmiZdm7G+IZQuPvTNsmfH3Aj4ie04kPijJfoVG0vfUiEaK/IKEJ6JeM66ZLKHr+5PCUIoLdvH
IsEUJLXhiiaxcm9X/+AbAF3fJtIUPclMiWckR2e31kGQ0cI1kRtP6eyWYo+XfHV2hK2gNCup6k2a
1ddh2Y+aq6Lvge6RnLOqau1e+HLYsaXYKK0SOcfZXRwcE+sELeERBFoTlBmhXZwV592UaMqyEG4T
sFalqkxdfTV2U6eOFAb6cBVKylA2TY2vqBIyYyRpt0+/Z/hWYtU4e5/SKVoWlSAi2TYN08qe8Zoj
cCGanTXkT5YOM53tSJ3vGmQZ038AgA+8pBgcSqSM64c34foTX77n2BwbWjywNOgIv8sc4qVmAz6q
u/t9SgffblluAsOaDEmd6gq8R56FN+nqeOJOyvIJoTMUdOHp+rEe8mRUAzCKC60L2XEMMWk7sDYI
3d7OJ4kjWLHDItRA77+T66Pz99CYaIJ4hVcgR7KOssEi08AB33CKs7xI/zC/0faI+SMwUUqKWYzU
Cy+4uqd5PA3IT+byoQ5bLrhQKIXg4rgQH5tJJ8338k/LnGRTNDeAyHSc3kbPlVSrsO8HdT1X4koW
eANcz3vXQOUrYIzKOOPq3gcPda+Y/rGzA0z1jK2lWW64wYm9Q3kPO3FJhSEyLy9GZ4UX8mjtWL2x
TPcnC77PG0ZqozOWCZ8XY1b6PahhDa9GY7DyETI6z3/V7BXX3bXhg7ysW4h1Vovh6jAfIgqYFURO
693Zt/M7LbigEQN5IndL7/8is8MMD2s4sN1+rffvru7RDnmFNE4liTwtf9UMTpvc2z/fPblWHc/d
PYtTw4qq6oAWaoouxW8fPD//UjQ5LQnTQi/FSC4S7m/klQNRtajZLnCaKDBad+dp3kTTUZtrhzoG
MOprEMx4r8GpOqtz0dc+8+QafPro7hbymSRKDR2Ldg7Ozg76fdmpgOHEOZ6aPQmfCEy65GVWzEuF
YZjfOHycAyoCrwd/7UQ25iUw0vzCtlQSma0NjUhyfom5hVx+T1cSHOb/Ay+sLk27JSk9Hbb+yOH8
cKGEsy6Pq88EoVN+AxtXEhbCdXs0QBDUMRV6MN5fdueeYJQSu85VGUUuOR7TDLGSzMRie909R2GC
FoDLPAL2mCYa5jwfGH5Io5UHek59YcHd/L04EFu2keyKqaaHurQ9OJxYXtFfD4fVnIV4ez/H4uZV
KBqB8GS+PBb29giqLvXG3G10wQB2e+O4kpAxsms3PHpBcw8NiqELyOA9apUnlTYd2tlXabcuGxQT
C5lJlyf2B6uclI0y9sbO2XqTXiAzLbwpuDSbF3/CC1Sgy98BfQ0pUtZbGSmMVNhhsfX53sJh8p53
/Y8MeH6l59IMUn/Mt47Da63OqtAsaVXOevcyIg3YOLmg0t3gLBpOwWpFexUQdKh61j5PwI1QQh/Z
9PAJF0FTHgBw40fGUpLeYQDqyRFXSNnQgw5L/Qx+PU4YlVSMb4FL07LShKTMbImXu0+yISEVyZsq
Izkqjx/7GKsrPu5bMonuEhE5FliI+RwcLRgB5YhyT8fkvZLdCcbmgoNqxYtGCtS4TqZljrPRK5b1
37bLlplHtIW9YTGlly+6YoJa+DPzOE8QarYRa6UztmfTtcpXhXms5A1Xc/EoJ/bnqxGiwtX6ghrv
BhvR+n/ILfGD7GdAlr9ksW9+Ien567TqJZkUknLYnOVegI6bvW53U3Rx54LQBtonaTmTrfzJqWGV
XeJ46v127UKtAmGj/CgKUZQb9nf2NMb0YcGHDiNU3T80RCABLKILbF29Kch24BBgzSZGzp7p1loF
cLH3HrnI4iKjLuJR4hk3rgAu97olxlo2t0qNb2kROAlT50rXHeTmuiH0WmTBnViuyF+B90quDC6Z
YRj144e8U7iqfA2hZLNYel04qrwEGBnaogJJ55dGNST0f40uVd3PS6aBNNfKSHhKNsi0ylM0u1aj
1q9LDrN+saSNNvZb5S7iRUPskh++7Clcpa7Vk3AwfR5+dCuzN1lM2s14R+sxsZgbvRUyem0hrT7i
hJFn33824uXZ6DOSNrcCIygMsHyFRJrP2IrwNqC9MC2XanJQHPB4+4Ay66rzd55VVcGKJi22yXeO
Mjd0auqOlVgCGXtiVlAQSkkEtGsG8hC/QC0dezsohNG+6lBtIWsFLXU38TUh3ZIAzG50g5JxnrG9
m7uPRB0FEAc6tPF8LtQ10kHr/x0VTONyy6Q779W1Bb+g36McA3XoVKoon8fWq0qR4Pia8SmmIu72
o+NNPu8qxe57rIXIFcsvKwFxGxg/Y6Pg6zfxa8KdE9zao9CR59goMmo7jc/AhJo1Y09L6Jj/KWDB
CjzU6p09r6y7ycp4g3r28sj24cUAbGwVFzI/pFvp3JQm1dhTf5ExvuX3RsVOGlCPWwCXJvtvygY5
SLG77NDC3BEMYnwVeSSzSClTBjr0l35bP78JgBxplx9XfLaMY1fCWczATI3YPxoNgzv1sreuD7V0
/6ZrtXzmowqrydXonHUIDW0eHuMWZp4eDEzxE+3T9+N5HEvcYKsQHGgsONUZ0aUaNTY6lF6EPKlD
rmtjJyIYr8bBQW1mPWsqDBki9AbD5UZHd0icUYLA3x96pgN96sWiE1iHPImdB93oGUS8B2E+NM1U
pRxX/hDnBeQFdkTyijRJ3jNj2GjEHyuRMiEohoSHtaolTnuxWD9IoniZ5UMFT06Q8YdbcY8QO0MY
7N4kdnCM
`protect end_protected
